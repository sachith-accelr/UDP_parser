// ************************************************************************************************************************
//
// Copyright(C) 2022 ACCELR
// All rights reserved.
//
// THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF
// ACCELER LOGIC (PVT) LTD, SRI LANKA.
//
// This copy of the Source Code is intended for ACCELR's internal use only and is
// intended for view by persons duly authorized by the management of ACCELR. No
// part of this file may be reproduced or distributed in any form or by any
// means without the written approval of the Management of ACCELR.
//
// ACCELR, Sri Lanka            https://accelr.lk
// No 175/95, John Rodrigo Mw,  info@accelr.net
// Katubedda, Sri Lanka         +94 77 3166850
//
// ************************************************************************************************************************
//
// PROJECT      :   40Gbps UDP Parser
// PRODUCT      :   NA
// FILE         :   UDP_NONBLOCKING_tb.sv
// AUTHOR       :   Sachith Rathnayake
// DESCRIPTION  :   Test Bench for UDP parser
//
// ************************************************************************************************************************
//
// REVISIONS:
//
//  Date           Developer               Description
//  -----------    --------------------    -----------
//  13-FEB-2023    Sachith Rathnayake      Creation
//
//
//*************************************************************************************************************************

`timescale 1ns/1ps

module UDP_NONBLOCKING_tb ();

    //---------------------------------------------------------------------------------------------------------------------
    // Global constant headers
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // parameter definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // localparam definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    localparam  ClOCK_PERIOD        =   6       ;
    localparam  BEAT_PERIOD         =   6       ;
    
    //---------------------------------------------------------------------------------------------------------------------
    // type definitions
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // I/O signals
    //---------------------------------------------------------------------------------------------------------------------
    
    logic   [255:0]         In_data         ;
    logic                   In_valid        ;
    logic                   Out_ready       ;
    logic                   clk             ;

    logic                   clkD            ;

    logic                   reset           ;
    logic   [255:0]         Out_data        ;
    logic                   Out_valid       ;
    logic                   In_ready        ;
    
    //---------------------------------------------------------------------------------------------------------------------
    // Internal signals
    //---------------------------------------------------------------------------------------------------------------------
    
    
    
    //---------------------------------------------------------------------------------------------------------------------
    // Implementation
    //---------------------------------------------------------------------------------------------------------------------
    
    UDP_NONBLOCKING udp (
            .In_data            (In_data  )     ,  
            .In_valid           (In_valid )     , 
            .Out_ready          (Out_ready)     ,
            .clk                (clk      )     ,      
            .reset              (reset    )     ,    
            .Out_data           (Out_data )     , 
            .Out_valid          (Out_valid)     ,
            .In_ready           (In_ready )         
    );
    
    initial begin
        clk         =   1'b0    ;
        forever begin
            #(ClOCK_PERIOD/2)   clk = ~clk      ;
        end
    end

    initial begin
        clkD        =   1'b0    ;
        forever begin
            #(BEAT_PERIOD/2)   clkD = ~clkD      ;
        end
    end

    initial begin
        
        @(posedge clk)  reset       =   1'b0    ;
        #1              reset       =   1'b1    ; 
        
        
        @(posedge clk)  Out_ready   =   1'b1    ;
       
        //-- First packet arravial--

        // while (!In_ready) ;
            //In_valid    <=      1'b1;
           if (In_ready) begin
               @(posedge clkD) In_valid = 1'b1;
                               In_data <= 256'h0034_0026_0006_0014_0040_0028_001D_0008_0030_002E_003D_0023_0001_0022_0022_0028 ;
               @(posedge clkD) In_data <= 256'h002F_001E_000C_001C_000D_0002_000C_000D_001E_0023_0021_001B_002D_0004_001E_0038 ;
               @(posedge clkD) In_data <= 256'h003C_001F_001D_001A_001D_0007_0023_003E_0001_0002_0014_0030_0025_000A_000B_0006 ;
               @(posedge clkD) In_data <= 256'h000C_0007_0021_0024_000C_0025_0006_0029_003E_003F_001C_0012_001B_000A_003D_0006 ;
               @(posedge clkD) In_data <= 256'h0035_000F_0017_0026_003D_0018_000D_0016_0003_0007_000D_000A_0014_0015_0026_0001 ;
               @(posedge clkD) In_data <= 256'h0040_0032_0019_0000_0034_0031_003C_002E_0015_0024_0026_002C_002A_003D_0021_0030 ;
               @(posedge clkD) In_data <= 256'h002C_000F_000B_0012_0027_0008_003A_0008_000B_0020_002C_002C_0013_0000_0022_0007 ;
               @(posedge clkD) In_data <= 256'h0025_0023_0026_0014_0001_0016_003D_0018_002B_0035_0017_0022_0012_0022_0015_0007 ;
               @(posedge clkD) In_data <= 256'h0041_0028_0031_0000_0039_0041_0022_0040_0011_0038_0036_0008_002D_000B_0028_000C ;
               @(posedge clkD) In_data <= 256'h0006_0017_001F_0032_001B_000F_0000_0031_0037_000A_0004_002D_000B_0007_0002_0021 ;
               @(posedge clkD) In_data <= 256'h0024_0024_001E_0027_0039_0032_0034_0034_0033_000A_0006_0025_002F_000E_000D_000E ;
               @(posedge clkD) In_data <= 256'h0020_001C_0006_0017_003C_0013_0018_0035_0035_0012_0004_0040_0038_0040_003B_000C ;
               @(posedge clkD) In_data <= 256'h0021_003A_0038_0001_001F_0041_0033_003D_003D_001D_000F_0034_001C_0025_0035_0026 ;
               @(posedge clkD) In_data <= 256'h002B_000B_002D_0005_0035_003F_002C_0007_0024_000E_002D_0011_0019_0041_001E_0037 ;
               @(posedge clkD) In_data <= 256'h0027_003D_003E_0037_0033_0028_0019_002A_0027_003C_0037_0000_0029_0001_000B_000E ;
               @(posedge clkD) In_data <= 256'h001A_0016_0026_0000_000E_000C_0008_0012_001D_0011_003A_0002_0039_0018_0038_0022 ;
               @(posedge clkD) In_data <= 256'h0027_0022_0005_001E_0010_0002_002F_0003_0002_0012_0022_000D_0030_0041_0037_0034 ;
               @(posedge clkD) In_data <= 256'h0015_000A_0010_0035_0024_002F_003B_0033_0005_0030_0022_001C_0035_0037_002B_000C ;
               @(posedge clkD) In_data <= 256'h0004_0013_0018_0024_002D_0006_0017_000C_0005_0024_002B_0013_002E_0025_0034_0021 ;
               @(posedge clkD) In_data <= 256'h003D_002A_0034_0001_000A_0011_003B_0038_002E_0028_0001_0016_0037_0009_002D_001A ;
               @(posedge clkD) In_data <= 256'h0034_000D_0016_002C_0040_001E_0016_003D_0003_0022_000D_0039_0036_000A_0017_0041 ;
               @(posedge clkD) In_data <= 256'h000D_0023_001D_003A_003A_0011_0007_001A_0011_0006_0024_0001_0039_002C_000F_0002 ;
               @(posedge clkD) In_data <= 256'h002E_0018_0015_001C_0016_0025_0009_0007_0006_0038_001C_003A_002A_002C_0008_002B ;
               @(posedge clkD) In_data <= 256'h003F_0032_0006_0035_0015_0040_0004_0031_0031_0002_002D_0032_0012_0021_0006_003B ;
               @(posedge clkD) In_data <= 256'h0005_002A_0032_0001_0018_000D_002F_0013_0020_0006_0021_001F_000C_001A_0034_0027 ;
               @(posedge clkD) In_data <= 256'h0028_0004_0016_0005_0005_003D_003E_001F_0021_000F_001C_002C_0001_002D_0015_001B ;
               @(posedge clkD) In_data <= 256'h0031_0041_0027_0025_000F_0041_000F_0015_0002_003D_0022_003C_001A_0013_0026_0028 ;
               @(posedge clkD) In_data <= 256'h0012_0006_0028_002E_0020_0017_0033_0020_0016_0007_003A_003E_003F_0040_003F_003F ;
               @(posedge clkD) In_data <= 256'h0012_000A_003A_0030_0028_002A_001C_0005_000C_000C_0034_0018_0021_000E_000A_001D ;
               @(posedge clkD) In_data <= 256'h0028_0016_0019_003E_0010_003C_0026_0012_0009_002D_0009_002D_0027_0014_0028_0007 ;
               @(posedge clkD) In_data <= 256'h000E_0016_0005_0031_0019_0010_0010_001B_000B_0041_0029_000D_0036_0027_0001_0016 ;
               @(posedge clkD) In_data <= 256'h003C_0028_0038_003E_0040_000A_0041_0030_0024_000D_001C_000E_002B_0020_0017_001B ;
               @(posedge clkD) In_data <= 256'h0017_001B_002E_0005_003E_0026_0012_000E_0033_0027_0002_002C_0006_002D_0008_0003 ;
               @(posedge clkD) In_data <= 256'h0005_002A_0019_0038_000A_0039_0003_0022_0034_000A_0000_000A_0027_001D_003C_002A ;
               @(posedge clkD) In_data <= 256'h002C_0025_000C_003A_0002_0022_0025_0022_000C_002D_0027_0032_0010_0018_0011_0018 ;
               @(posedge clkD) In_data <= 256'h0017_0004_0034_0034_0021_000E_0014_003A_0000_0038_0025_000E_0026_003D_0026_002E ;
               @(posedge clkD) In_data <= 256'h003F_0017_003D_0008_003C_001E_0016_0007_000A_0031_0005_000C_003A_0035_002C_0034 ;
               @(posedge clkD) In_data <= 256'h001C_0034_000F_0025_0039_001C_0002_0031_0038_003C_0031_0007_0012_003C_001E_0010 ;
               @(posedge clkD) In_data <= 256'h000D_0025_000B_0010_0008_0014_003F_001B_0001_0025_0041_003A_0000_0018_0035_0028 ;
               @(posedge clkD) In_data <= 256'h0036_0000_001F_002B_001D_000C_0016_0009_002C_0016_001B_0004_0005_000A_0015_0008 ;
               @(posedge clkD) In_data <= 256'h001F_0014_0015_0009_0035_0002_0004_0027_0037_0020_0004_0029_001F_0028_0040_002E ;
               @(posedge clkD) In_data <= 256'h0037_0026_0026_000C_0035_0021_0002_002A_0005_002C_0028_003F_001F_0000_0000_000E ;
               @(posedge clkD) In_data <= 256'h0032_0017_002B_0005_000D_0030_0016_001E_0019_003C_0017_0001_0009_0006_0023_002A ;
               @(posedge clkD) In_data <= 256'h0038_0016_0031_0017_003F_000F_0039_000E_0014_0001_003E_0004_0000_0014_000C_003E ;
               @(posedge clkD) In_data <= 256'h001B_0004_001C_0014_0035_0011_001E_0039_0005_000A_0015_002A_0021_0013_003F_002D ;
               @(posedge clkD) In_data <= 256'h001F_0016_0021_0000_002C_000C_0023_0033_002D_000B_003C_002C_0006_0041_0036_0029 ;
               @(posedge clkD) In_data <= 256'h001B_0008_001D_0017_000B_003C_0038_0011_0014_0009_0028_0010_0027_000C_003D_0041 ;
               @(posedge clkD) In_data <= 256'h0032_0014_0005_0027_0003_0006_0015_0027_002C_0022_0020_0015_0021_0009_0032_0036 ;
               @(posedge clkD) In_data <= 256'h000B_003C_0013_000C_0003_0035_002C_0022_001A_0017_0041_0004_0033_001C_0006_0018 ;
               @(posedge clkD) In_data <= 256'h0003_0034_002F_0018_001C_0025_0010_002F_0014_003C_0018_003C_0007_001A_002C_0012 ;
               @(posedge clkD) In_data <= 256'h003F_0011_0041_0001_0001_001B_001F_001C_001C_001F_0013_002C_001F_003A_002F_0003 ;
               @(posedge clkD) In_data <= 256'h0037_0031_0004_001C_0016_0004_0035_0024_001C_0034_002D_000B_002B_0035_003D_0017 ;
               @(posedge clkD) In_data <= 256'h0026_001C_0026_000D_0007_0030_0014_0038_001A_003F_0016_000B_0030_002A_0011_0037 ;
               @(posedge clkD) In_data <= 256'h000A_0008_0038_0026_001E_0023_0018_003A_003A_0010_0039_0020_0029_0002_0009_0039 ;
               @(posedge clkD) In_data <= 256'h002A_003A_002D_001D_000C_0030_002A_003A_0021_0031_001D_0039_0018_0008_0024_0021 ;
               @(posedge clkD) In_data <= 256'h001B_0031_000D_0005_000B_0004_001C_003C_0034_0025_001E_0021_0011_0030_0033_000C ;
               @(posedge clkD) In_data <= 256'h001B_0000_000F_001E_0002_0020_0033_000F_002A_002A_003F_0041_0013_0035_001B_0029 ;
               @(posedge clkD) In_data <= 256'h0000_0007_0028_0004_0035_0028_0029_001E_001A_002F_000E_0006_003B_003D_0041_0038 ;
               @(posedge clkD) In_data <= 256'h001F_0001_002D_0028_002C_0001_0022_003D_0040_002D_002D_000A_000A_0007_0034_0014 ;
               @(posedge clkD) In_data <= 256'h002F_0015_001F_000C_0032_000A_001E_0027_000E_001A_0020_0020_0032_000B_0020_0034 ;
               @(posedge clkD) In_data <= 256'h0010_0015_0013_0038_0038_0020_0004_000B_002E_0041_0000_0019_0031_0028_0041_0037 ;
               @(posedge clkD) In_data <= 256'h001C_001B_003B_000B_000E_0017_0010_000E_0003_0012_000D_0037_0035_0015_0020_003B ;
               @(posedge clkD) In_data <= 256'h0019_001C_0013_000F_0016_003C_002F_003A_0000_0000_0000_0000_0000_0000_0000_0000 ;    
           end
           

      // @(posedge clkD)Out_ready   <=   1'b1 ; 
       // end of packet

      // @(posedge clkD)
       //  In_valid    <=      1'b1;
       //output is ready
       

      // while (!In_ready) ;

          //2nd

            if (In_ready) begin
                @(posedge clkD) In_valid    <=      1'b1;

                                In_data = 256'h0002_0030_0009_002D_0031_000F_0008_001E_0012_000A_003C_0026_0032_001D_001F_0034 ;
                @(posedge clkD) In_data = 256'h000D_0027_002E_0037_002A_0001_000C_002B_0009_002E_0012_0009_002C_001B_0000_0019 ;
                @(posedge clkD) In_data = 256'h0020_0029_003B_0030_0030_002A_001B_0024_0009_0023_001B_0018_0011_003C_0011_0039 ;
                @(posedge clkD) In_data = 256'h002E_0002_000D_000D_0020_000B_001D_003E_0023_0033_0004_0030_002D_0008_0039_0037 ;
                @(posedge clkD) In_data = 256'h0040_0011_0021_0005_002A_0010_0008_001D_0009_0030_000A_0003_0037_0027_0030_002A ;
                @(posedge clkD) In_data = 256'h0032_0001_0012_003F_0015_0029_0011_0025_0017_002A_0012_0000_0032_0039_003F_0038 ;
                @(posedge clkD) In_data = 256'h000F_000E_0007_0018_0039_0027_000A_0008_0036_0032_0016_0036_000E_0008_001F_0035 ;
                @(posedge clkD) In_data = 256'h002F_0013_0007_003F_0038_0020_001D_0036_0027_0015_0019_0005_0006_0014_0001_000E ;
                @(posedge clkD) In_data = 256'h0007_0000_0031_001D_0001_000A_002C_0020_003C_003D_0023_0026_002A_000F_0010_0007 ;
                @(posedge clkD) In_data = 256'h0020_000A_0006_0006_000A_001C_0008_0028_002F_0016_0040_0033_0028_0017_0011_002E ;
                @(posedge clkD) In_data = 256'h0022_0021_0039_0025_001F_003F_000D_0036_003A_0027_003B_000A_0017_0040_003C_0038 ;
                @(posedge clkD) In_data = 256'h0002_0022_000B_0007_003C_000F_0024_000A_0037_0037_002B_0036_0023_0016_001A_001C ;
                @(posedge clkD) In_data = 256'h000A_000F_001F_0023_001C_003A_0039_002A_0027_0024_002B_0012_0032_0008_0039_0021 ;
                @(posedge clkD) In_data = 256'h003B_0009_0032_0038_0023_0021_002F_0010_0005_0020_000A_0019_003A_0040_0019_0006 ;
                @(posedge clkD) In_data = 256'h0011_0023_002E_0016_002C_0015_0013_001F_0040_0004_0034_000C_0020_0041_0035_0009 ;
                @(posedge clkD) In_data = 256'h0035_0016_003F_000A_0013_002E_0026_003D_0003_003F_0036_003A_0016_0002_003B_002B ;
                @(posedge clkD) In_data = 256'h002C_000E_0010_000D_0002_002C_000D_0019_0005_0037_0008_002B_0003_0004_0001_0002 ;
                @(posedge clkD) In_data = 256'h002A_003A_0034_0035_0024_0002_0011_000D_0017_0007_0002_0016_0011_002A_0010_003D ;
                @(posedge clkD) In_data = 256'h0021_0011_001B_002E_0028_0036_000A_0041_0018_0022_0031_0041_0040_000F_000B_003C ;
                @(posedge clkD) In_data = 256'h0038_0018_003E_0027_0011_003C_0001_002A_002B_0016_0013_001D_0041_002B_001B_0036 ;
                @(posedge clkD) In_data = 256'h0041_002F_0009_0034_0031_002B_0033_003E_0000_0027_0018_000E_000B_0018_000B_0011 ;
                @(posedge clkD) In_data = 256'h002C_003C_0017_0005_0013_0007_0009_0003_0004_0021_0038_0009_001D_000E_000B_0033 ;
                @(posedge clkD) In_data = 256'h0008_0015_0017_0007_0016_0032_002D_0012_0021_0015_0001_0028_0020_0020_0032_0032 ;
                @(posedge clkD) In_data = 256'h003D_0018_0016_0030_0008_002A_0025_000A_0022_0033_002C_0038_002E_0009_0023_001D ;
                @(posedge clkD) In_data = 256'h001C_003D_0037_0030_0028_001A_003B_0024_0010_0030_0033_001D_0017_0019_0008_0000 ;
                @(posedge clkD) In_data = 256'h003E_0016_0006_003F_0010_000D_000E_001A_0023_0016_002C_0001_000F_0009_0016_003D ;
                @(posedge clkD) In_data = 256'h0019_001D_0011_0019_000D_000A_0015_0030_0028_0022_0000_0033_0003_0041_003F_0018 ;
                @(posedge clkD) In_data = 256'h0031_0010_001D_0029_0002_0025_0029_0003_001F_003F_0007_001E_0000_0027_000E_0038 ;
                @(posedge clkD) In_data = 256'h0013_0016_003F_0018_0031_003D_001E_0020_003F_0020_0017_0022_000E_002A_001D_002A ;
                @(posedge clkD) In_data = 256'h0014_0005_001D_0035_001B_0005_000B_0000_0032_0024_0016_001E_0027_0035_000B_0003 ;
                @(posedge clkD) In_data = 256'h0008_0029_003E_0027_0036_0036_0016_0040_0032_0041_0028_0000_0007_002D_0019_001B ;
                @(posedge clkD) In_data = 256'h0022_000C_0030_0002_000D_0026_0019_0009_0005_000A_0041_0033_001E_0035_0022_0028 ;
                @(posedge clkD) In_data = 256'h003B_0019_003E_001C_0021_002D_002E_001B_001D_002B_001D_001B_0002_000D_0032_003A ;
                @(posedge clkD) In_data = 256'h0026_002C_0023_0018_0041_0000_0021_000D_0000_0037_0018_0006_0035_002E_0021_0040 ;
                @(posedge clkD) In_data = 256'h003F_002F_0008_0037_0033_0002_0037_0013_003F_0034_0021_000E_0027_0015_001B_0007 ;
                @(posedge clkD) In_data = 256'h002B_000E_0015_003D_0036_002F_002D_0031_001D_002A_0028_002D_003D_003B_0030_0000 ;
                @(posedge clkD) In_data = 256'h0028_002A_000C_0038_001B_0015_0007_001A_0031_000D_001B_000B_0009_0024_003F_002D ;
                @(posedge clkD) In_data = 256'h001A_0031_002B_0017_0001_0037_0010_003B_0001_0024_000F_001C_0013_0001_003D_000A ;
                @(posedge clkD) In_data = 256'h0003_001C_002F_0031_0000_0003_0016_003C_002C_003C_0026_000E_0029_001C_0030_0027 ;
                @(posedge clkD) In_data = 256'h000F_0008_0013_0020_0040_0001_003D_001E_0027_002E_0002_0027_002F_0029_0004_0027 ;
                @(posedge clkD) In_data = 256'h0033_002C_0029_0014_000D_0034_002E_0023_0007_0039_0004_0041_001C_0008_0001_000A ;
                @(posedge clkD) In_data = 256'h0040_0038_000A_0013_0034_0021_0020_0041_000C_001E_002B_0038_0036_0013_0021_001C ;
                @(posedge clkD) In_data = 256'h0027_001E_001A_001C_0037_0000_0021_0029_0026_0014_0000_000E_0008_003B_0039_0034 ;
                @(posedge clkD) In_data = 256'h0039_0026_003C_001D_0007_0026_0031_003D_0011_0027_0033_0013_0004_0014_0023_0011 ;
                @(posedge clkD) In_data = 256'h0025_0028_0029_001F_0000_0010_0028_0036_0005_0023_0014_0003_0003_0019_003D_003B ;
                @(posedge clkD) In_data = 256'h0038_0040_0022_002B_0033_0000_0038_0007_0005_001C_0018_0034_0029_0032_0040_0019 ;
                @(posedge clkD) In_data = 256'h0022_0017_0038_0025_0008_003E_0040_0027_0004_0036_0037_0020_002E_0020_0016_003A ;
                @(posedge clkD) In_data = 256'h0021_0015_002E_001C_001B_0008_0001_0016_0024_0038_000A_0029_0032_0041_0037_000F ;
                @(posedge clkD) In_data = 256'h0039_0003_000B_000A_0011_0036_0003_0004_0002_001E_0018_0010_003F_0022_0003_0036 ;
                @(posedge clkD) In_data = 256'h000D_0003_0039_000B_003B_0018_001A_001B_001C_002B_002A_0034_003B_0020_001B_0024 ;
                @(posedge clkD) In_data = 256'h0036_0038_0016_0011_0009_002A_0020_000B_0038_000C_000C_0035_0035_0019_002B_0030 ;
                @(posedge clkD) In_data = 256'h0035_003B_0011_0024_002F_0036_001A_0041_0021_0022_000B_0009_0039_002B_0011_003E ;
                @(posedge clkD) In_data = 256'h002E_0016_0009_0000_003A_0038_001E_0005_0019_000E_002D_0005_002B_0031_0022_0031 ;
                @(posedge clkD) In_data = 256'h000B_0034_001F_001F_0038_0028_0036_0040_0011_001A_0018_0014_0041_003F_0030_000C ;
                @(posedge clkD) In_data = 256'h003F_0025_0013_0030_0005_0006_0034_0007_0028_0001_0006_0022_0002_0038_001F_0039 ;
                @(posedge clkD) In_data = 256'h0034_000C_0026_0037_0035_0020_0021_001D_003B_0013_0013_0004_0001_0018_0008_0035 ;
                @(posedge clkD) In_data = 256'h0007_003B_0012_000A_0031_0010_003A_0019_0025_0026_001F_0027_0027_0031_0037_0010 ;
                @(posedge clkD) In_data = 256'h0034_0008_0005_0035_0010_0036_000B_001B_0022_001F_003D_000B_0012_0005_0005_0036 ;
                @(posedge clkD) In_data = 256'h001A_000A_0035_0027_001A_000E_0011_0011_0002_0037_0014_003B_0014_002C_000A_0012 ;
                @(posedge clkD) In_data = 256'h0011_001C_0005_0024_0011_0012_001C_001E_0025_0033_003F_003E_003B_0013_0009_0038 ;
                @(posedge clkD) In_data = 256'h0036_0034_0033_003C_0021_0021_0009_000B_002F_001C_003C_003C_0040_0023_0023_0040 ;
                @(posedge clkD) In_data = 256'h0014_000F_000F_003C_0029_0018_0027_0009_0027_0027_0012_002A_001E_0003_0035_001E ;
                @(posedge clkD) In_data = 256'h0015_002B_002C_0018_000F_002D_0032_0027_0000_0000_0000_0000_0000_0000_0000_0000 ;
            end



        // @(posedge clkD) Out_ready   =   1'b1 ;
        
        // end of packet
        // @(posedge clkD)

        //In_valid    <=      1'b1;
        //output is ready
        
        // while (!In_ready) ;

            //3rd

           if (In_ready) begin
                @(posedge clkD) In_valid    <=      1'b1;

                                In_data = 256'h0015_0031_003D_0017_0032_0028_0001_0012_0009_0018_001A_0012_002B_0004_0028_0004 ;
                @(posedge clkD) In_data = 256'h000D_0037_0018_000E_0013_0001_000C_0011_0016_0009_0027_0040_0012_003C_0002_0012 ;
                @(posedge clkD) In_data = 256'h0022_000D_002F_001D_0010_0010_0009_003F_003E_0016_0017_0004_003C_0029_002A_0026 ;
                @(posedge clkD) In_data = 256'h0036_0016_0029_0018_0017_0038_0034_0040_0025_0030_000B_0008_0007_0017_001E_0006 ;
                @(posedge clkD) In_data = 256'h0030_0024_0026_003D_0003_0040_002C_001E_0007_0008_0025_001D_003D_002B_000D_001F ;
                @(posedge clkD) In_data = 256'h0008_001D_0035_001E_002C_0039_0023_0022_000B_003B_0017_0020_0009_0018_001F_0012 ;
                @(posedge clkD) In_data = 256'h0005_002F_0017_000C_0016_002D_0040_0029_0036_0009_0007_0027_0030_0013_0038_002B ;
                @(posedge clkD) In_data = 256'h0036_0009_0021_003F_003A_0010_0026_0018_0014_0040_0017_0024_000A_0003_0015_0034 ;
                @(posedge clkD) In_data = 256'h0020_0039_0025_003F_0002_0005_0026_002E_000C_002C_0015_002D_0006_0041_0038_0016 ;
                @(posedge clkD) In_data = 256'h0009_0038_0020_0017_001A_0011_000B_0014_0026_0020_0007_0011_002B_003E_0002_0036 ;
                @(posedge clkD) In_data = 256'h0003_0041_0040_0024_000F_0038_001C_0019_003D_0005_001E_003B_001A_001F_003E_002D ;
                @(posedge clkD) In_data = 256'h000C_0003_0033_0037_0039_001F_0022_002C_003E_0002_001F_0018_003D_0027_0019_0039 ;
                @(posedge clkD) In_data = 256'h0030_0014_0024_0012_001F_0007_0019_003E_000D_0038_0004_003E_001E_0009_0007_000C ;
                @(posedge clkD) In_data = 256'h001B_002E_001E_000C_0006_0030_003E_0023_0029_001B_000C_002D_001C_0001_0022_0016 ;
                @(posedge clkD) In_data = 256'h000F_003A_0009_003A_0023_0003_001B_0035_0015_0035_002B_0000_0035_0033_0029_003A ;
                @(posedge clkD) In_data = 256'h0013_0019_002A_0019_0033_001E_003C_0030_0015_002C_003E_0006_001A_0010_0008_000B ;
                @(posedge clkD) In_data = 256'h0000_002F_0021_0026_001A_0008_003F_0010_003F_0028_0040_0000_0005_000A_0024_0008 ;
                @(posedge clkD) In_data = 256'h0003_0017_0029_001D_0018_0003_0030_0022_001C_0032_0035_002E_0036_0034_0040_0002 ;
                @(posedge clkD) In_data = 256'h002D_003F_0019_000D_001F_0006_0004_0003_000B_0036_0033_0013_0003_002E_000B_002C ;
                @(posedge clkD) In_data = 256'h0037_003E_002C_0019_001E_000B_0040_0017_003D_0036_001C_0014_000E_002E_0019_002A ;
                @(posedge clkD) In_data = 256'h0018_0009_003F_0017_003B_0041_000D_003D_0016_0017_002C_002F_0030_0020_0036_000B ;
                @(posedge clkD) In_data = 256'h001B_001E_001C_0003_0027_003C_0021_0005_0035_0000_0018_001A_0015_0012_000F_0030 ;
                @(posedge clkD) In_data = 256'h002A_0006_0032_001C_0013_001D_0012_0013_0034_002E_0031_0015_003E_0030_0019_0037 ;
                @(posedge clkD) In_data = 256'h002C_0023_0035_001C_003A_003B_002C_001F_001D_002C_0010_003D_0008_001B_003B_003A ;
                @(posedge clkD) In_data = 256'h000C_0002_0006_0019_001F_0041_000F_0018_0007_000B_0015_0001_0003_0014_0027_001F ;
                @(posedge clkD) In_data = 256'h0016_0005_0034_0028_001D_0028_002B_000F_002C_002C_0022_0012_0025_0010_0007_002B ;
                @(posedge clkD) In_data = 256'h002D_003A_001E_001F_0001_001F_001E_0001_0028_003C_0037_0035_0018_000F_0032_0005 ;
                @(posedge clkD) In_data = 256'h000B_0035_000C_0034_002B_000C_0025_0028_001A_0011_002E_0033_0034_0006_001E_0034 ;
                @(posedge clkD) In_data = 256'h0007_001E_001A_0014_000F_0000_0020_0014_0001_0028_0010_003E_0004_000B_0010_003E ;
                @(posedge clkD) In_data = 256'h000B_0012_0040_0005_0006_0018_0033_0037_002C_000E_0017_0037_0031_000E_003D_0009 ;
                @(posedge clkD) In_data = 256'h0028_0011_003A_0008_0031_001C_0025_0013_0000_001B_003A_003E_0006_002F_0001_0029 ;
                @(posedge clkD) In_data = 256'h0018_0012_002D_000A_000F_0029_003B_0018_000E_001A_0038_002E_001A_0027_002C_0028 ;
                @(posedge clkD) In_data = 256'h003B_002F_0003_002C_0032_0017_0016_0006_0002_002D_001A_003B_000F_0020_0032_000B ;
                @(posedge clkD) In_data = 256'h002C_0012_001B_001D_0006_0023_0015_0011_001E_0033_003A_0023_0041_002B_0002_0012 ;
                @(posedge clkD) In_data = 256'h0004_0031_0026_0001_001A_0001_0017_003F_003A_001A_0036_000C_0012_001A_0039_003E ;
                @(posedge clkD) In_data = 256'h0035_002E_0027_0017_001D_0010_003B_001E_0021_0017_0014_001E_002B_000D_0009_0014 ;
                @(posedge clkD) In_data = 256'h0029_0034_0016_0008_0026_000C_0004_003A_003C_000D_001D_000C_0019_003B_002B_0021 ;
                @(posedge clkD) In_data = 256'h000F_0030_000B_0000_0017_0005_0019_002F_0005_0023_0037_003E_0016_0036_002C_0026 ;
                @(posedge clkD) In_data = 256'h000A_0014_003C_0003_0009_002C_0027_0027_000A_0018_003E_0026_003A_002B_002F_0035 ;
                @(posedge clkD) In_data = 256'h001F_0025_001C_0040_0001_0021_002F_0005_002B_0041_0017_0021_000D_003B_0030_003B ;
                @(posedge clkD) In_data = 256'h0001_003D_0012_0019_0033_0024_0029_0026_002B_001A_0004_000B_002A_003A_000A_0017 ;
                @(posedge clkD) In_data = 256'h000A_000E_001F_000D_0000_0010_0018_0030_0007_002F_0027_0036_0010_0020_003C_0027 ;
                @(posedge clkD) In_data = 256'h0039_000E_0013_003A_0039_002D_0025_000E_001F_003B_0022_003D_003C_000D_0000_0030 ;
                @(posedge clkD) In_data = 256'h0007_0010_0035_0000_001E_000E_001F_0033_0028_0031_002A_0025_0027_0031_0035_000D ;
                @(posedge clkD) In_data = 256'h003A_000F_000C_0029_002E_0008_000B_001E_0007_0028_0040_002F_000A_003B_0028_0023 ;
                @(posedge clkD) In_data = 256'h0033_0009_0039_001D_0032_0003_002F_0014_0040_0036_002E_0021_002E_002F_002A_001F ;
                @(posedge clkD) In_data = 256'h003B_0011_0027_003E_0030_0032_002E_0018_0037_0015_0028_0022_0023_001F_003B_0004 ;
                @(posedge clkD) In_data = 256'h0016_0006_0028_0019_0025_0010_0009_0036_0026_002F_0010_0033_0003_002F_001F_003B ;
                @(posedge clkD) In_data = 256'h0014_0030_0001_002D_001C_0015_0000_0020_0040_002B_0012_0013_003B_0000_0000_0019 ;
                @(posedge clkD) In_data = 256'h0008_0038_0004_0041_001A_001C_000E_0026_0036_000D_0000_0025_003D_0016_0039_0024 ;
                @(posedge clkD) In_data = 256'h002F_001E_0002_0016_0004_0016_0002_000A_001D_0000_0005_0008_0030_0007_0004_000C ;
                @(posedge clkD) In_data = 256'h002C_0002_001F_0012_002D_002B_0036_003E_0021_0021_000C_0041_0033_0014_001C_000B ;
                @(posedge clkD) In_data = 256'h001C_0037_002B_0035_002A_0033_000A_0004_0037_0016_0010_0019_0010_0016_002F_000F ;
                @(posedge clkD) In_data = 256'h0033_002D_0028_0038_0039_0035_002C_002E_001A_000C_000E_0018_0038_0010_0022_0031 ;
                @(posedge clkD) In_data = 256'h0032_002E_0007_0011_0010_003B_0029_0010_002B_003D_003F_003C_000B_0032_0012_0028 ;
                @(posedge clkD) In_data = 256'h0000_0022_0032_0008_0008_0029_003A_0020_0008_0033_0008_000F_0025_0022_001A_000F ;
                @(posedge clkD) In_data = 256'h003C_0005_0028_001F_0001_0032_0032_0026_0041_000A_0023_0038_0001_000C_0008_003F ;
                @(posedge clkD) In_data = 256'h001D_0003_0034_0031_002B_0017_0030_0038_002B_0002_001F_001F_0016_0021_0035_0009 ;
                @(posedge clkD) In_data = 256'h0040_0001_0025_0006_0001_0007_000C_0008_0037_0020_0036_003E_0035_0010_0037_0022 ;
                @(posedge clkD) In_data = 256'h0026_0024_0026_0014_003F_002B_003B_003B_003E_000D_0034_003C_002E_0039_0008_002F ;
                @(posedge clkD) In_data = 256'h001B_002F_003E_0040_0026_001E_0037_0025_000B_002F_0004_002A_0031_0007_001A_0019 ;
                @(posedge clkD) In_data = 256'h0006_0021_002F_003A_0009_0034_002C_0005_0020_0007_0039_0026_0032_0037_002C_001F ;
                @(posedge clkD) In_data = 256'h0036_0031_0022_0032_0005_0022_000E_000D_0000_0000_0000_0000_0000_0000_0000_0000 ;
           end
        
        // @(posedge clkD) Out_ready   =   1'b1 ;
        
        // end of packet
        // @(posedge clkD)
        //In_valid    <=      1'b1;
        //output is ready

        // while (!In_ready) ;
            //3rd

                // 4th

            if (In_ready) begin
                @(posedge clkD) In_valid    <=      1'b1;

                                In_data = 256'h0029_002B_0021_0006_0015_0036_0008_0011_0005_0018_0002_0014_0024_0041_000A_003B;
                @(posedge clkD) In_data = 256'h0027_000D_0005_0025_0010_0002_000C_0016_003A_0040_002D_0018_0001_000A_0039_000A;
                @(posedge clkD) In_data = 256'h0017_003A_000B_0041_000C_000B_003A_0002_0019_0032_002C_003A_0032_0020_000E_000D;
                @(posedge clkD) In_data = 256'h0013_000D_0039_0014_0001_000F_001E_0001_0024_002D_0001_001A_0027_000C_0015_0004;
                @(posedge clkD) In_data = 256'h0029_003C_0011_001E_003E_0031_002F_0002_002F_001E_0023_0015_002A_0033_0008_001A;
                @(posedge clkD) In_data = 256'h0039_0007_0019_000B_001B_0034_0001_0023_002A_0006_0004_0036_0034_0010_0013_003E;
                @(posedge clkD) In_data = 256'h0039_000C_0034_0041_0001_000E_000F_0014_000E_003F_000B_0026_0033_000D_0027_001E;
                @(posedge clkD) In_data = 256'h0037_0033_0021_001E_002C_0024_0016_0008_000C_0039_0039_0020_0022_0032_002E_0036;
                @(posedge clkD) In_data = 256'h0015_0022_0039_0021_001D_0022_0030_0029_0017_002F_0030_0012_0036_0029_0016_0017;
                @(posedge clkD) In_data = 256'h0005_0006_002F_0041_003E_002D_0009_000E_0030_0039_001D_0026_0016_0005_0019_000D;
                @(posedge clkD) In_data = 256'h0003_0011_0029_0010_0027_0002_000A_002D_0017_0017_001A_0009_001F_0014_0041_001F;
                @(posedge clkD) In_data = 256'h0028_0025_0009_0041_0021_002C_002A_0040_0003_0001_0037_0029_0014_0018_000E_0036;
                @(posedge clkD) In_data = 256'h0009_0014_000E_0020_0032_0034_003D_000C_001C_0000_0014_0035_0040_0036_000B_0004;
                @(posedge clkD) In_data = 256'h0022_0031_000A_001B_0026_0011_0005_0040_002A_0037_0031_0015_0035_0010_0025_0000;
                @(posedge clkD) In_data = 256'h0017_002B_001E_001F_002F_0009_003F_0024_0016_0014_0041_0024_0021_0029_0008_0005;
                @(posedge clkD) In_data = 256'h003F_002C_0009_000A_0024_000F_003C_002D_0033_000C_0013_0034_0033_0017_0017_0003;
                @(posedge clkD) In_data = 256'h0039_000B_0011_002A_0014_003B_0033_001A_0028_0002_001A_0012_0000_0036_001C_0011;
                @(posedge clkD) In_data = 256'h0009_0013_000C_0031_0041_000B_0013_0014_0006_001C_0031_001E_0038_0013_0028_0023;
                @(posedge clkD) In_data = 256'h0015_0016_001D_0017_003B_0013_0037_0031_0015_0025_002B_0034_0031_0035_0025_0016;
                @(posedge clkD) In_data = 256'h002E_0015_003A_0011_0010_003C_0023_000A_003C_000C_0041_0038_0014_0025_0021_0033;
                @(posedge clkD) In_data = 256'h001B_002A_0036_003C_000C_0031_0011_0025_0014_001E_0026_002B_0028_0017_002F_001B;
                @(posedge clkD) In_data = 256'h0041_0038_0012_0041_000B_0012_001C_0028_003A_0021_000F_0019_0037_003C_002B_0020;
                @(posedge clkD) In_data = 256'h002F_0027_0017_0037_0028_0027_000D_0009_0003_0023_0005_0015_0031_0039_0023_0028;
                @(posedge clkD) In_data = 256'h0025_000D_0038_0031_0031_0038_0040_0001_0035_0014_003A_0014_0040_0024_0019_0016;
                @(posedge clkD) In_data = 256'h0009_000A_0008_0028_0019_003D_0034_0000_001F_003C_0011_0033_002C_0004_0039_0036;
                @(posedge clkD) In_data = 256'h001C_003E_0015_002F_0019_003A_0037_0002_002B_000F_002E_0018_000B_0023_002D_003B;
                @(posedge clkD) In_data = 256'h0023_0025_0033_000C_0022_0011_0030_002A_0000_002D_002F_0009_0009_002D_0032_003B;
                @(posedge clkD) In_data = 256'h0041_0037_0037_003D_0033_0001_0012_001D_003E_0025_0007_0020_0040_0016_000E_000C;
                @(posedge clkD) In_data = 256'h003F_000A_0018_0041_002A_0010_003E_0036_001A_0032_0011_0013_001B_001F_001F_003A;
                @(posedge clkD) In_data = 256'h003A_0012_0030_0005_000F_002B_0020_0030_0029_0021_0036_0025_001F_001E_000A_001A;
                @(posedge clkD) In_data = 256'h000D_003A_0031_000C_0004_0019_001C_0032_0023_0034_003B_0012_0004_0026_0027_003F;
                @(posedge clkD) In_data = 256'h0023_002C_0030_0015_001B_002F_0040_0019_0002_002E_0025_001E_002D_0041_000F_0026;
                @(posedge clkD) In_data = 256'h0041_0040_0037_001A_0028_002E_0040_001F_003E_0000_000C_0034_0003_0010_0003_0000;
                @(posedge clkD) In_data = 256'h0032_0034_002F_0001_0008_0022_002E_001C_0024_000E_002D_001B_0006_0034_0036_003F;
                @(posedge clkD) In_data = 256'h0033_0021_000D_0038_0008_002D_003F_003A_0016_000E_0034_0033_0010_001A_0032_0036;
                @(posedge clkD) In_data = 256'h002B_0020_0021_0033_000B_0005_000A_0007_0016_0015_000C_0030_0015_0002_0006_002B;
                @(posedge clkD) In_data = 256'h0004_0005_003C_0034_0020_0014_0018_0000_0030_001D_002A_0037_003D_0041_0008_003B;
                @(posedge clkD) In_data = 256'h0004_000E_001E_0007_002B_000B_0003_001E_0028_0011_0015_0019_002F_002B_0041_000C;
                @(posedge clkD) In_data = 256'h0039_0002_001F_0040_0040_0022_0035_0002_0011_0029_002A_0015_002D_003B_0028_0029;
                @(posedge clkD) In_data = 256'h0009_0009_0030_0024_0014_002C_0032_002D_001B_001B_000E_0029_003B_0001_0029_0033;
                @(posedge clkD) In_data = 256'h0039_0000_0022_0007_0021_0001_001A_0036_0005_003E_0004_001E_0021_003B_0013_0034;
                @(posedge clkD) In_data = 256'h0037_0014_0028_003A_0014_0028_0031_003C_002E_002A_0016_002B_003B_0020_0041_001A;
                @(posedge clkD) In_data = 256'h0024_0027_0029_0021_000F_0011_0028_000D_000F_0031_001A_0001_000F_0021_0015_003A;
                @(posedge clkD) In_data = 256'h0035_0013_0033_0004_002D_0013_0041_0012_003E_003C_0020_0027_001A_0000_0033_0023;
                @(posedge clkD) In_data = 256'h000E_0025_0037_002C_0020_0020_0029_0007_0005_003B_001E_0004_0002_002D_0015_0000;
                @(posedge clkD) In_data = 256'h001A_001E_0004_001B_002E_000B_0021_002C_0036_0009_001E_0025_001E_0003_0036_0018;
                @(posedge clkD) In_data = 256'h0034_002B_0037_002A_0028_001B_002C_0034_003A_0034_0026_001C_002A_0012_0022_0024;
                @(posedge clkD) In_data = 256'h003D_0019_0007_000D_0029_003D_001D_0010_000E_0001_000D_0030_002D_0025_0001_001B;
                @(posedge clkD) In_data = 256'h0021_002A_0007_0027_0035_0018_0029_0010_0021_0039_001C_0019_003F_0029_003A_003E;
                @(posedge clkD) In_data = 256'h0034_001C_0012_0017_0011_0030_0023_0020_0031_0037_000D_003D_0028_002D_0010_0004;
                @(posedge clkD) In_data = 256'h0022_002D_002E_000E_002A_000B_003A_003D_001C_0038_0002_003B_000A_0013_003D_003C;
                @(posedge clkD) In_data = 256'h001E_0040_0023_001C_0016_003F_0028_0034_0029_0021_0031_0040_001F_0015_003C_000E;
                @(posedge clkD) In_data = 256'h0014_0018_0018_0017_0005_002A_0024_000A_0039_003E_003E_002D_0002_0004_0026_0001;
                @(posedge clkD) In_data = 256'h0033_0016_0009_0006_0019_0034_0029_0002_001A_0040_0031_003D_002D_0004_0033_000E;
                @(posedge clkD) In_data = 256'h003D_0017_000F_0001_0011_0017_001C_0010_0031_000C_0027_003D_0021_0032_0007_0033;
                @(posedge clkD) In_data = 256'h0009_003F_0037_0025_002D_0041_0023_0030_0011_0011_001F_002D_0031_0038_000C_0000;
                @(posedge clkD) In_data = 256'h0041_0004_0005_003F_0039_0017_0037_002B_0040_003E_0011_0014_0008_000A_0014_0030;
                @(posedge clkD) In_data = 256'h0041_000E_0028_0014_0016_0035_0009_001E_0036_000E_0003_0025_001C_0034_0022_002E;
                @(posedge clkD) In_data = 256'h0022_001A_0038_003B_0019_002E_0027_0012_0036_0032_0015_0001_0010_0003_0010_0016;
                @(posedge clkD) In_data = 256'h0029_000B_0041_0024_0003_0040_0018_0008_0016_0003_0023_002D_0028_0036_002B_0026;
                @(posedge clkD) In_data = 256'h0005_003C_002C_0018_002E_0004_0015_001D_0036_0008_000C_0035_0037_001D_001C_003B;
                @(posedge clkD) In_data = 256'h0013_003F_0009_000C_0006_003D_0015_0031_003A_001B_0036_003F_001E_0030_0022_0006;
                @(posedge clkD) In_data = 256'h0005_003F_0016_0015_0012_0033_0024_0013_0000_0000_0000_0000_0000_0000_0000_0000;
            end
            // end of packet
            // @(posedge clkD)
            //output is ready
        

        // @(posedge clkD) Out_ready   =   1'b1 ;

        // while (!In_ready)  ;


            // 5th

        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;

                            In_data = 256'h000B_0032_001D_003D_0008_0005_0021_0024_0037_0027_002B_000B_003C_001F_001C_0022;
            @(posedge clkD) In_data = 256'h0036_0041_002C_002D_0012_0002_000C_003D_0021_0030_0022_000D_0028_0001_0027_0000;
            @(posedge clkD) In_data = 256'h0006_002B_0040_003C_000D_003E_0027_000E_0031_0032_0010_001D_0004_0011_000C_0036;
            @(posedge clkD) In_data = 256'h0018_001C_002D_000B_003C_0009_002F_003D_0029_0003_0022_0010_0003_0035_0012_002C;
            @(posedge clkD) In_data = 256'h0006_001D_0025_0015_003B_000C_0015_000B_0000_003E_0035_0029_0022_003C_003E_0032;
            @(posedge clkD) In_data = 256'h0014_001E_0003_0003_0004_0003_0034_0028_001E_0039_0020_0023_0009_002A_0039_0022;
            @(posedge clkD) In_data = 256'h0040_0007_0002_0039_0009_002E_0025_0004_001C_0018_0014_002A_0040_000A_001D_0037;
            @(posedge clkD) In_data = 256'h0038_001A_001E_0008_0020_001F_002E_0012_0012_0035_0034_0010_0021_0039_0019_001B;
            @(posedge clkD) In_data = 256'h0002_002A_0027_002A_000B_0003_000B_0008_0005_003F_001D_0037_000D_0035_0035_002B;
            @(posedge clkD) In_data = 256'h003B_0003_0020_003D_003A_003B_0038_000C_001F_002D_0010_002B_003E_0010_0018_003B;
            @(posedge clkD) In_data = 256'h0008_0025_0016_0021_0007_0031_0011_0013_003A_0005_0013_000B_001D_0012_001A_0010;
            @(posedge clkD) In_data = 256'h0005_003A_001F_0011_000C_0008_0034_003F_0032_0019_003C_0039_0027_003A_001F_0021;
            @(posedge clkD) In_data = 256'h001A_001F_0000_0040_0038_0012_003F_0019_0020_0032_0013_0035_0012_0014_0001_0035;
            @(posedge clkD) In_data = 256'h0010_000F_0005_003F_002A_001F_0016_0038_000D_0012_0009_002D_0015_0012_0016_0005;
            @(posedge clkD) In_data = 256'h0025_0013_0010_003B_003E_0023_0035_000C_0029_0011_002A_000C_0032_0035_0011_003E;
            @(posedge clkD) In_data = 256'h0023_0001_0019_0004_000A_0019_0012_003D_0001_0004_001B_0005_0002_0036_0006_003A;
            @(posedge clkD) In_data = 256'h0035_000B_0010_0026_0026_0040_0033_0041_0011_0040_000A_0013_002C_0032_0000_0029;
            @(posedge clkD) In_data = 256'h0021_002B_0028_000A_0002_003D_003C_0011_000E_001B_001C_0012_003E_0041_0005_0009;
            @(posedge clkD) In_data = 256'h002C_001A_001D_003F_002E_0032_002F_0022_0038_0036_0007_0021_0016_0034_0030_0022;
            @(posedge clkD) In_data = 256'h0019_002C_003A_0013_002D_002C_0016_000D_0002_000B_0021_0005_0014_0027_0026_001B;
            @(posedge clkD) In_data = 256'h002C_0018_0011_0023_002D_001B_002A_000F_0004_002D_000D_0023_002A_001D_000C_0001;
            @(posedge clkD) In_data = 256'h0015_0041_0040_001E_0012_0025_003C_001E_0031_003D_0003_0034_0016_003A_001B_002A;
            @(posedge clkD) In_data = 256'h0032_003A_0019_0021_0001_0027_0040_003C_0012_001E_0032_000B_0032_0011_0013_003E;
            @(posedge clkD) In_data = 256'h000A_0036_002D_0036_0025_003F_0032_0017_002D_0037_0040_000D_002D_0038_002D_0021;
            @(posedge clkD) In_data = 256'h003D_002B_001F_0001_0020_002F_001E_0032_0018_0033_0031_0032_0041_002D_0007_0006;
            @(posedge clkD) In_data = 256'h003F_0036_0006_001B_000F_0008_0029_0004_0013_001C_000A_0033_0028_0015_0035_0034;
            @(posedge clkD) In_data = 256'h001A_0022_0023_0041_000C_001D_0034_0023_0002_0035_0023_000C_000D_0025_0015_000F;
            @(posedge clkD) In_data = 256'h0021_0020_0033_0028_0008_001A_0039_0034_002D_002F_003A_0006_0015_0009_001A_003A;
            @(posedge clkD) In_data = 256'h001D_0028_003A_0035_000A_0033_001C_0041_0021_0023_0009_003F_000E_0041_0022_000B;
            @(posedge clkD) In_data = 256'h0024_002E_0015_0019_0039_0039_003D_003B_0028_001A_003F_0027_001D_0003_001B_0004;
            @(posedge clkD) In_data = 256'h0022_002E_0006_001B_001E_0025_002C_0017_003B_0038_0037_0034_003B_0035_000E_002B;
            @(posedge clkD) In_data = 256'h0022_0013_0001_0038_002D_0030_001D_0035_0007_0022_0025_0023_0009_001E_0013_0035;
            @(posedge clkD) In_data = 256'h0021_002C_0004_0015_0023_0003_0014_001D_0017_003A_0017_0037_0019_0008_000F_0035;
            @(posedge clkD) In_data = 256'h0014_000A_0009_0015_000F_002A_0037_000B_0006_0004_003E_003D_003E_003E_001E_0037;
            @(posedge clkD) In_data = 256'h0018_0023_0022_002E_0037_0015_0018_002C_0006_0003_000D_000D_0030_0006_001E_0020;
            @(posedge clkD) In_data = 256'h0038_0025_0009_002A_003B_001D_0017_0003_0039_0031_001E_0002_000A_0025_0024_003C;
            @(posedge clkD) In_data = 256'h0033_0034_002F_002B_0039_003A_0035_001D_0020_002F_002A_0027_0034_0033_003B_0003;
            @(posedge clkD) In_data = 256'h0036_001D_0017_0005_001A_0012_002A_001A_002D_003C_003E_0019_0001_0006_000F_0029;
            @(posedge clkD) In_data = 256'h0016_0028_0017_0014_0032_000F_0025_0015_0018_0013_0030_0019_001A_0035_0025_0000;
            @(posedge clkD) In_data = 256'h0005_0008_0026_002E_002D_0022_0035_0027_000B_003D_0027_0029_002B_002D_002E_0038;
            @(posedge clkD) In_data = 256'h0025_000A_003F_0007_0006_003E_000C_001B_0032_0019_0004_0029_0015_0037_003B_003A;
            @(posedge clkD) In_data = 256'h0000_0030_002A_003A_001C_0033_0041_0035_000A_002C_0031_003B_0038_0036_0025_0030;
            @(posedge clkD) In_data = 256'h0039_000B_0005_001B_0031_0002_0038_0028_0008_000E_003A_001E_0039_0025_002D_000C;
            @(posedge clkD) In_data = 256'h0033_000F_0025_003D_0016_0001_000E_0005_0023_0029_001A_0010_0012_000E_0003_002E;
            @(posedge clkD) In_data = 256'h0018_0001_0034_002B_0014_0012_000C_0018_0014_002F_0010_000D_0028_0041_0005_000D;
            @(posedge clkD) In_data = 256'h003A_001D_0028_001F_0039_001E_002C_0035_0014_0034_0017_003C_000F_0018_003D_001F;
            @(posedge clkD) In_data = 256'h003B_0022_001F_001C_0004_001D_0036_0003_0021_0008_0002_000C_0031_000B_002D_0019;
            @(posedge clkD) In_data = 256'h0034_0003_0029_0020_0002_0008_0015_002E_0019_002D_001A_000A_0020_0022_001E_0010;
            @(posedge clkD) In_data = 256'h0014_003E_0003_0005_000F_0009_0035_0025_0012_0041_0004_0009_0023_0021_002A_0032;
            @(posedge clkD) In_data = 256'h000B_0008_001F_0020_0039_0022_003D_0005_0018_001A_001F_0004_0020_003B_0037_003F;
            @(posedge clkD) In_data = 256'h003C_0023_0024_0004_0030_0021_001D_0039_0014_003C_0000_0032_0038_0014_0006_002A;
            @(posedge clkD) In_data = 256'h001E_0001_002C_003C_0025_0024_0022_0006_000A_0029_0036_002E_001A_001D_0022_0009;
            @(posedge clkD) In_data = 256'h001B_003A_0036_001A_0041_0010_002A_0016_000D_003F_0005_0026_000F_0024_0005_000D;
            @(posedge clkD) In_data = 256'h0013_0029_0003_0022_001D_0031_0031_0038_002E_0012_0037_0011_0040_0010_001A_0030;
            @(posedge clkD) In_data = 256'h0015_0004_0014_0019_0021_0032_000A_0011_0002_003D_003F_0026_0032_0008_0039_0014;
            @(posedge clkD) In_data = 256'h0012_0009_003A_0021_000B_0020_0026_0023_001B_0006_0016_003D_0041_000D_0012_0021;
            @(posedge clkD) In_data = 256'h0017_000D_003F_0035_0024_0010_0029_0000_0003_001D_003A_0037_0007_0011_0000_003A;
            @(posedge clkD) In_data = 256'h0018_0004_0034_0023_001D_0004_002E_0003_002D_002E_0040_002C_0040_0020_000F_003A;
            @(posedge clkD) In_data = 256'h0011_0015_000B_0022_002C_0029_0003_000E_0003_003B_0022_0015_0009_000C_0016_0010;
            @(posedge clkD) In_data = 256'h0033_002A_002D_0034_0016_0020_0003_001A_000E_0010_0034_0039_001B_002D_0029_001A;
            @(posedge clkD) In_data = 256'h0039_0008_002E_003E_0001_0032_0009_000A_0010_0001_0007_0026_0026_0039_002C_0020;
            @(posedge clkD) In_data = 256'h0025_0002_0040_001D_0016_000C_0004_0017_002F_0034_0041_0001_0005_000B_0032_0011;
            @(posedge clkD) In_data = 256'h0005_003E_0003_0027_0005_003E_001B_002F_0000_0000_0000_0000_0000_0000_0000_0000;
            
        end    
            // end of packet
            // @(posedge clkD)
            //output is ready
        

        // @(posedge clkD) Out_ready   =   1'b1 ;

        // while (!In_ready)  ;

        // 6th
        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;

                            In_data = 256'h002A_0008_0004_001A_0009_002D_0009_0015_0008_000F_0010_001B_0041_000E_002D_0012 ;
            @(posedge clkD) In_data = 256'h0037_0026_0018_002A_0038_0001_000C_002B_0021_0021_001A_0024_001F_003D_0041_0012 ;
            @(posedge clkD) In_data = 256'h001F_003C_0019_0005_0039_000D_0041_0011_0040_002C_0022_0025_0021_0027_0010_0008 ;
            @(posedge clkD) In_data = 256'h0035_0017_000B_0019_0024_0032_0016_0012_0006_0017_003E_0041_0005_0002_000D_0020 ;
            @(posedge clkD) In_data = 256'h001D_0029_000A_0010_0009_0025_0006_0026_0032_0025_0010_0015_001F_0019_0035_0035 ;
            @(posedge clkD) In_data = 256'h001A_0017_0020_0009_0040_0040_0017_003F_0030_0019_0030_001F_0022_0036_000C_0038 ;
            @(posedge clkD) In_data = 256'h0027_0033_0002_0019_000E_0013_000E_001F_0019_001D_0009_0017_003E_001F_002F_001E ;
            @(posedge clkD) In_data = 256'h0029_0020_0011_0017_0037_0004_002D_0020_001C_0038_0027_001F_0011_0030_0031_0038 ;
            @(posedge clkD) In_data = 256'h0041_0004_0028_002C_0013_003C_0036_001F_0001_001D_0014_000B_0015_002C_0029_0025 ;
            @(posedge clkD) In_data = 256'h0036_000D_0037_0008_0028_000A_003D_001E_002D_002F_000C_0008_003A_003C_0020_0017 ;
            @(posedge clkD) In_data = 256'h0002_001F_001E_001B_0003_001B_0016_0025_0010_0034_000B_002E_000F_0035_001F_0026 ;
            @(posedge clkD) In_data = 256'h0039_000D_0012_0016_000D_002F_0020_0022_0004_0008_0018_003B_002C_003D_0021_0035 ;
            @(posedge clkD) In_data = 256'h002A_002E_0005_000A_003D_0007_0039_002A_002B_0022_0024_0039_0016_002D_0041_0033 ;
            @(posedge clkD) In_data = 256'h0010_0025_0034_000E_0007_0041_0033_001E_0035_001C_002A_0021_0017_0011_0018_0017 ;
            @(posedge clkD) In_data = 256'h0021_0013_0001_0023_0025_003C_0030_0011_0006_0017_002E_000F_0011_0016_003C_0018 ;
            @(posedge clkD) In_data = 256'h0022_0028_0032_0034_000B_0009_002B_002C_001B_0035_0038_0031_001C_0002_0012_0040 ;
            @(posedge clkD) In_data = 256'h002F_001A_000D_0019_0000_001B_0014_003C_0028_0021_0028_0002_0034_003C_001A_0006 ;
            @(posedge clkD) In_data = 256'h0034_0005_0029_000C_002A_0031_0030_0004_0018_002B_0014_000E_0012_001F_001F_0019 ;
            @(posedge clkD) In_data = 256'h001B_0024_000E_003C_0018_0023_0035_002B_0018_0027_0001_001A_0014_0027_0026_0026 ;
            @(posedge clkD) In_data = 256'h0001_0041_0007_003E_0010_000E_0013_001C_0017_0013_0031_0005_000B_0009_0012_0021 ;
            @(posedge clkD) In_data = 256'h002C_0020_0011_000D_0003_0029_003C_002C_003B_003D_002F_000C_002C_0013_001D_003B ;
            @(posedge clkD) In_data = 256'h003D_0008_0020_0018_0040_0025_0008_0034_001D_0014_0016_0030_0022_002E_000F_003B ;
            @(posedge clkD) In_data = 256'h001E_0013_0005_0038_001F_0035_002E_000D_0031_0009_0031_0029_0007_0002_001D_0033 ;
            @(posedge clkD) In_data = 256'h0025_0021_0007_0039_003B_0017_002C_0029_0024_0016_0031_000E_0010_002C_0032_0016 ;
            @(posedge clkD) In_data = 256'h0009_003D_0019_0023_0031_0000_0002_003A_0033_002C_0001_0021_0012_0006_003B_0006 ;
            @(posedge clkD) In_data = 256'h0025_0016_003F_000A_0004_003A_0010_0005_0018_0001_0041_0028_003C_0009_003E_0005 ;
            @(posedge clkD) In_data = 256'h0008_002C_001D_0005_0012_0038_0009_0029_0035_003B_000C_0020_001C_0008_000E_002B ;
            @(posedge clkD) In_data = 256'h0007_0004_001C_001E_001E_001A_0035_0009_0033_0041_0016_0010_0028_0034_0018_0012 ;
            @(posedge clkD) In_data = 256'h0000_002C_0021_0012_0027_0022_000A_0015_0010_001C_000E_003A_0014_002E_0040_0037 ;
            @(posedge clkD) In_data = 256'h0025_000D_0008_0013_0028_002B_0030_0006_0021_000D_0021_001C_0000_002D_000A_0023 ;
            @(posedge clkD) In_data = 256'h000C_0001_0019_0033_0034_003C_0004_002E_001D_0025_0039_0003_003F_0027_0041_0021 ;
            @(posedge clkD) In_data = 256'h0027_0031_0027_003A_003C_0016_0008_000F_003C_0028_0013_0016_0028_002C_0010_0007 ;
            @(posedge clkD) In_data = 256'h002C_002A_0015_0009_0022_002F_001A_0002_0032_0021_0038_0032_0001_0039_0002_0033 ;
            @(posedge clkD) In_data = 256'h001D_003E_0003_0013_0031_0023_001F_0009_0021_002A_0024_002F_0010_000A_000D_0024 ;
            @(posedge clkD) In_data = 256'h0033_0035_0023_001D_0021_0021_0037_0012_003E_0016_002C_000B_0012_0003_0002_0003 ;
            @(posedge clkD) In_data = 256'h0029_0013_003C_002F_0006_0030_002C_0005_001F_0039_0035_002A_0023_0005_0006_003E ;
            @(posedge clkD) In_data = 256'h002D_000A_002F_0028_003A_000B_0025_003B_002E_0038_0030_0002_0009_0035_0030_0023 ;
            @(posedge clkD) In_data = 256'h002E_002C_002D_0012_0001_0012_002A_0032_001D_0001_0031_0018_003B_0025_0010_0020 ;
            @(posedge clkD) In_data = 256'h0019_000C_0024_0001_000A_0036_001F_000D_002D_0030_001F_0016_0025_0004_0036_0004 ;
            @(posedge clkD) In_data = 256'h003F_000F_002D_0040_0014_0034_003F_0014_000B_0002_0019_0020_001D_0033_000E_001D ;
            @(posedge clkD) In_data = 256'h001D_002D_0003_0026_0023_0018_001A_002A_0028_0028_0004_002E_0014_0011_0023_003D ;
            @(posedge clkD) In_data = 256'h000C_003B_0001_000D_000D_003A_0032_002B_0034_003F_003D_0026_0022_0024_000A_0026 ;
            @(posedge clkD) In_data = 256'h0038_0000_000B_0040_0005_0024_0015_002E_0006_001E_0033_003D_000D_0004_003A_003E ;
            @(posedge clkD) In_data = 256'h0004_001C_001C_0005_0016_000D_0001_0029_0025_0009_000B_0040_0011_000C_003D_0001 ;
            @(posedge clkD) In_data = 256'h0026_0025_0031_0033_0020_0038_0007_0020_0000_000B_0011_002E_0037_003D_0002_0007 ;
            @(posedge clkD) In_data = 256'h003B_0025_0018_003A_0001_000A_0033_003F_0034_0026_0029_0015_001B_002D_0006_0012 ;
            @(posedge clkD) In_data = 256'h0006_0027_0018_0009_0012_000F_0000_0031_0021_002C_003D_0031_000E_002D_0004_0024 ;
            @(posedge clkD) In_data = 256'h000D_0022_003C_0022_0037_000E_0013_001D_002A_0029_0013_0020_000F_001F_0031_0006 ;
            @(posedge clkD) In_data = 256'h0026_0005_000B_0017_0022_0014_001E_0024_001D_001D_0004_0029_0020_0004_0025_0004 ;
            @(posedge clkD) In_data = 256'h0035_001A_0017_0022_0005_002E_001E_0000_001B_0000_000E_0019_0011_001B_0025_0018 ;
            @(posedge clkD) In_data = 256'h003B_0014_0036_0022_0007_0020_0021_0019_001C_001D_003F_0016_001B_0020_002A_000F ;
            @(posedge clkD) In_data = 256'h002D_0041_0041_001F_0020_000C_0018_000F_001E_0035_002B_0020_003C_0019_0018_003C ;
            @(posedge clkD) In_data = 256'h0040_0028_002F_0007_001A_0022_001B_0031_001C_002B_001F_0037_0018_0024_003B_0007 ;
            @(posedge clkD) In_data = 256'h0024_0010_000D_0011_003E_0036_0015_0023_001F_003D_0010_001F_0032_0005_0011_000F ;
            @(posedge clkD) In_data = 256'h001D_0028_0018_0017_0027_003F_002D_000A_0018_001C_0034_002C_0033_003B_003A_002D ;
            @(posedge clkD) In_data = 256'h002C_0000_003C_003E_001C_0031_002D_0004_000E_0034_0038_0000_0039_0031_0017_001B ;
            @(posedge clkD) In_data = 256'h0015_0017_0009_0027_0034_0007_001E_0019_0021_0029_000E_0008_0037_0022_003B_0001 ;
            @(posedge clkD) In_data = 256'h0006_0005_0007_003D_002F_0038_000A_0015_0007_0027_003A_0012_0004_0005_0017_003D ;
            @(posedge clkD) In_data = 256'h002C_0014_0039_0018_0013_0005_0030_0033_002E_0014_0019_0002_0009_001E_000B_003E ;
            @(posedge clkD) In_data = 256'h0014_001D_0000_000F_0030_0039_0035_0014_0001_000D_0022_0011_0014_0008_002B_0019 ;
            @(posedge clkD) In_data = 256'h0034_0038_0025_0019_0040_002C_0033_0041_003C_003D_0018_0015_0020_0041_0018_002E ;
            @(posedge clkD) In_data = 256'h0031_0031_0027_0006_0036_0005_001C_0018_001B_0012_001E_001B_003E_0018_0005_0001 ;
            @(posedge clkD) In_data = 256'h0027_002F_000E_0028_0002_001B_0015_000B_0000_0000_0000_0000_0000_0000_0000_0000 ;
        end    
            // end of packet
            // @(posedge clkD)
            //output is ready
        

        // @(posedge clkD) Out_ready   =   1'b1 ; 
        
        // while (!In_ready)  ;

        // 7th
        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;

                            In_data = 256'h002E_003C_0002_003C_0014_0009_0035_0009_002D_0016_001F_003A_0031_001A_0028_001A ;
            @(posedge clkD) In_data = 256'h002F_0040_0035_003E_0026_0002_000C_0006_0019_002D_0028_0039_0033_0013_002A_0034 ;
            @(posedge clkD) In_data = 256'h003B_003B_003A_0027_0013_002A_0037_0029_0037_0009_0011_0012_000D_0027_0037_000E ;
            @(posedge clkD) In_data = 256'h000F_000E_0001_001E_003F_0030_0018_0001_002E_001B_0014_002F_0004_0026_0015_0030 ;
            @(posedge clkD) In_data = 256'h0036_003C_001F_0002_0006_0013_0034_000B_0001_003F_000F_0033_002B_002E_001E_003D ;
            @(posedge clkD) In_data = 256'h0004_0013_0008_0030_0018_0028_0011_003A_002B_0023_0019_0034_0003_001F_0017_0020 ;
            @(posedge clkD) In_data = 256'h0032_000C_003B_000A_001D_0037_001E_0015_002C_0031_0017_0038_0002_003C_0022_0020 ;
            @(posedge clkD) In_data = 256'h002A_0027_0038_000F_001E_0024_0021_0023_003F_000D_0034_002D_002A_001E_0026_0035 ;
            @(posedge clkD) In_data = 256'h003E_001F_0004_0011_0002_002D_0020_002D_0034_000C_0006_0037_000E_0031_0026_002E ;
            @(posedge clkD) In_data = 256'h0003_0028_0023_0013_003C_000F_0005_0036_000B_0007_002F_0001_0014_0008_0026_0000 ;
            @(posedge clkD) In_data = 256'h0041_0003_0018_0022_0035_0027_002D_0016_001B_002B_0011_0032_0016_0021_0010_0018 ;
            @(posedge clkD) In_data = 256'h0040_000E_0025_0039_003A_001E_003B_0040_0013_0026_002E_0033_0007_0010_000A_0035 ;
            @(posedge clkD) In_data = 256'h0025_000C_0003_0025_000C_0026_0025_0012_0011_0000_000C_000F_0029_0036_0036_001A ;
            @(posedge clkD) In_data = 256'h0028_0024_003A_0037_003C_0041_0038_000C_0021_000B_0029_0020_0035_0037_0034_003C ;
            @(posedge clkD) In_data = 256'h0020_003F_0029_0005_0026_0011_0020_0020_001A_001D_0024_002A_003C_0039_002F_0032 ;
            @(posedge clkD) In_data = 256'h0002_001B_0032_0015_0035_002D_0031_0015_000B_001A_0040_0011_0024_0011_0007_0015 ;
            @(posedge clkD) In_data = 256'h002F_000A_0004_0031_0035_001C_001A_0026_002C_0008_001C_0020_001E_003F_0030_0016 ;
            @(posedge clkD) In_data = 256'h0026_0023_000F_001C_0028_000F_0000_0014_001C_0008_0035_0025_0007_0025_0020_002B ;
            @(posedge clkD) In_data = 256'h0010_003E_0002_0007_0010_0008_0022_003A_0027_0039_0039_0028_0015_001B_002D_0010 ;
            @(posedge clkD) In_data = 256'h000E_000C_0005_0037_0023_003B_0007_0022_0021_001A_001B_003F_0008_001C_0034_001B ;
            @(posedge clkD) In_data = 256'h0007_0014_0013_0034_0023_0026_0023_0005_003E_0014_000D_000E_000A_0032_0023_0015 ;
            @(posedge clkD) In_data = 256'h000F_0000_0035_001F_001C_002E_000B_0039_002B_0003_001F_0003_0030_001E_0016_0028 ;
            @(posedge clkD) In_data = 256'h002E_001D_000A_002C_000C_001D_0010_002E_0030_0029_0039_0038_0022_002B_0031_001D ;
            @(posedge clkD) In_data = 256'h003D_0038_0009_0004_001D_0013_002D_0027_0017_0036_0002_001A_0028_0035_001F_0035 ;
            @(posedge clkD) In_data = 256'h0003_0022_0017_0009_002C_0018_0021_0014_0030_0037_0000_0022_0000_0022_0006_001D ;
            @(posedge clkD) In_data = 256'h0000_0004_0003_002F_003D_0018_0033_0012_002F_0020_0000_001F_003B_0020_003F_0037 ;
            @(posedge clkD) In_data = 256'h0040_0020_0025_003A_0028_0004_0017_0039_0035_0004_0003_0028_0032_0025_0034_0039 ;
            @(posedge clkD) In_data = 256'h0038_0014_0005_0033_0014_000D_0037_0007_0004_001E_0000_0037_0002_0001_002D_0035 ;
            @(posedge clkD) In_data = 256'h0001_0015_0020_001D_0039_002C_0009_0012_0031_0024_0040_0022_0031_000E_002F_003C ;
            @(posedge clkD) In_data = 256'h000D_0022_0006_0013_0023_0013_0031_0003_003E_001A_0039_0006_0033_003A_0019_002C ;
            @(posedge clkD) In_data = 256'h002B_0024_000F_0003_0023_002B_0016_0013_0035_0038_0000_0023_0030_002E_001D_003B ;
            @(posedge clkD) In_data = 256'h0023_0038_0018_000A_003C_002B_0041_0018_0005_003D_0009_0022_0038_003B_000F_0000 ;
            @(posedge clkD) In_data = 256'h001A_0002_0001_0006_002D_0040_0019_000A_0008_000C_003F_0008_0014_0004_0004_0024 ;
            @(posedge clkD) In_data = 256'h003E_0039_000D_0017_0012_0030_001C_001D_0035_000B_0009_000E_001C_001B_003A_0031 ;
            @(posedge clkD) In_data = 256'h0006_0010_0008_0033_0030_0013_0028_0006_0016_002D_001E_0006_0018_0041_002C_002B ;
            @(posedge clkD) In_data = 256'h002C_0025_002C_0017_0006_000E_0007_003C_0005_0035_002C_002C_003B_0017_0015_000E ;
            @(posedge clkD) In_data = 256'h0025_0026_0038_002C_0027_0019_003D_0010_0032_0002_001D_0040_003A_0007_0007_0021 ;
            @(posedge clkD) In_data = 256'h000E_003B_0014_002A_001B_0009_001C_0004_0003_003B_0016_0019_0007_0029_0015_002E ;
            @(posedge clkD) In_data = 256'h0021_0023_002D_002E_0021_0016_0018_0021_0027_0014_0038_0030_0019_0023_0000_0002 ;
            @(posedge clkD) In_data = 256'h0032_000E_0029_0019_0032_000B_001A_000A_0001_0005_001E_001F_0039_000A_0039_003C ;
            @(posedge clkD) In_data = 256'h002B_0035_0030_001F_0039_002C_002A_0025_001D_002F_0004_0023_0008_000A_0017_003F ;
            @(posedge clkD) In_data = 256'h0028_0007_003E_003E_0009_0039_0016_0034_000E_0009_0021_0004_0011_0009_002B_000A ;
            @(posedge clkD) In_data = 256'h000B_0022_0036_0002_0033_0016_002A_0027_0026_002D_003F_000B_0019_002E_001A_0041 ;
            @(posedge clkD) In_data = 256'h0021_0030_0031_0019_001F_0000_0014_001F_0033_0021_0026_0007_000C_002A_000E_0000 ;
            @(posedge clkD) In_data = 256'h0034_0033_0032_001F_0016_000F_0037_0037_0028_0005_0011_0002_0018_001C_0032_0028 ;
            @(posedge clkD) In_data = 256'h0001_0008_003F_0022_003D_0001_0018_001E_003B_0003_0023_000B_0041_002D_0012_002A ;
            @(posedge clkD) In_data = 256'h001A_0032_003F_0030_001C_002A_0029_0017_003F_001D_003D_0008_003F_0000_0009_0008 ;
            @(posedge clkD) In_data = 256'h0004_0029_000D_0029_0036_0018_0024_001A_0020_0021_003E_0026_0021_0010_0020_000D ;
            @(posedge clkD) In_data = 256'h0032_0016_003F_001A_0029_0015_0040_0034_000A_001D_0023_000B_003B_002B_0028_003A ;
            @(posedge clkD) In_data = 256'h0008_0038_0018_0012_003B_0031_0039_000D_0040_0008_001E_0037_0037_0037_0009_0032 ;
            @(posedge clkD) In_data = 256'h003B_003F_000C_0023_0007_0015_001F_003A_0004_0036_0018_0022_000D_0041_001B_0038 ;
            @(posedge clkD) In_data = 256'h001C_0041_0002_0002_0019_003E_0012_000B_0027_003E_001C_003E_0003_0002_0034_0014 ;
            @(posedge clkD) In_data = 256'h0009_0002_000B_0020_0011_0013_0004_001D_0020_0007_0041_001C_0012_0000_0027_001C ;
            @(posedge clkD) In_data = 256'h000C_000E_0016_001B_0004_003C_003A_0004_002C_0030_002E_0037_000E_0008_001F_001A ;
            @(posedge clkD) In_data = 256'h0035_002D_0035_001B_0039_0002_0014_000F_0007_003A_0031_0036_002E_0006_0039_002A ;
            @(posedge clkD) In_data = 256'h0036_0021_003C_0038_003C_0004_000A_0007_0026_003F_001B_0033_0036_0014_0027_0038 ;
            @(posedge clkD) In_data = 256'h002E_001D_0037_0026_003B_0006_001F_002C_000F_000B_003E_003B_0023_0002_0019_000D ;
            @(posedge clkD) In_data = 256'h0040_0033_0034_000B_000A_0026_0041_000F_0028_0029_0008_0017_000F_000B_0000_002F ;
            @(posedge clkD) In_data = 256'h000E_0005_0020_003B_0000_001A_0036_000A_001A_003A_001C_001D_0038_002E_003A_0003 ;
            @(posedge clkD) In_data = 256'h002C_0036_0022_0023_0022_0037_0011_0039_0022_0024_0036_0011_0013_0041_0025_0040 ;
            @(posedge clkD) In_data = 256'h0032_0033_0037_001B_001C_002E_0037_001F_000B_0007_003F_001B_0010_001C_001B_0039 ;
            @(posedge clkD) In_data = 256'h001F_0004_003E_002B_0028_0012_000F_0028_0014_001B_0021_0030_002F_0025_0008_0024 ;
            @(posedge clkD) In_data = 256'h003A_001D_0012_0034_0033_0028_0019_0034_0000_0000_0000_0000_0000_0000_0000_0000 ;
        end   
        // end of packet
        // @(posedge clkD)
        //output is ready
        

        // @(posedge clkD) Out_ready   =   1'b1 ;   

        // while (!In_ready)  ;

            // 8th
        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;

                            In_data = 256'h0023_0003_0004_0037_001F_0005_0014_003F_000E_002D_0009_003F_0017_0006_0009_0015;
            @(posedge clkD) In_data = 256'h0001_002F_001D_0022_0017_0002_000C_003F_0035_001F_0016_0038_0002_0019_0005_0036;
            @(posedge clkD) In_data = 256'h003B_0036_001E_0025_000C_000C_0025_0005_0041_0020_0015_0014_003A_003D_0014_000A;
            @(posedge clkD) In_data = 256'h0024_001F_001F_0026_0029_0037_0041_0021_0000_0035_000F_0002_0006_0004_000D_0023;
            @(posedge clkD) In_data = 256'h0012_002D_0038_0013_003F_0039_0008_0013_0021_001D_0011_000F_003A_0008_0020_0033;
            @(posedge clkD) In_data = 256'h0026_002A_0023_003A_002E_0014_000C_0012_0034_0020_0015_0006_002E_0002_0000_000F;
            @(posedge clkD) In_data = 256'h001A_003A_000F_0012_0010_0005_003E_0032_0009_000B_002A_0009_0030_0018_0003_0034;
            @(posedge clkD) In_data = 256'h0007_0023_0027_0033_003A_0034_002F_0038_002B_0031_0013_0041_000E_002B_0005_0017;
            @(posedge clkD) In_data = 256'h0032_002B_0005_0009_0021_0034_001D_0021_0036_0004_0041_0039_0002_0037_0003_0014;
            @(posedge clkD) In_data = 256'h0015_001C_000B_001D_0035_0037_0006_0036_001A_0035_000F_000A_0029_000B_0020_001F;
            @(posedge clkD) In_data = 256'h0006_002E_001B_003B_0010_003E_0000_002B_0021_0014_0008_0019_0040_0024_003B_003E;
            @(posedge clkD) In_data = 256'h0018_0035_0038_003B_0019_0001_0019_003F_0009_0008_0015_003E_000C_002C_0028_003A;
            @(posedge clkD) In_data = 256'h0022_0039_000A_0041_000F_000B_0002_0025_003D_0021_0001_0025_0024_0025_000B_0007;
            @(posedge clkD) In_data = 256'h0009_0022_0008_0023_000E_0035_001B_0026_0011_0038_0013_0024_0031_0015_0025_0029;
            @(posedge clkD) In_data = 256'h002E_003C_0024_001B_0037_0038_0031_0041_0031_0040_001A_0024_002B_0021_0018_0008;
            @(posedge clkD) In_data = 256'h0032_0019_002D_0023_001E_003F_003E_0012_0033_0022_0015_0029_0011_000D_0014_000C;
            @(posedge clkD) In_data = 256'h003D_002A_000C_0023_0024_0016_0007_0039_001C_000B_0018_003D_003A_000D_0000_002B;
            @(posedge clkD) In_data = 256'h003E_0038_0009_0002_000A_0025_0026_0009_001C_002F_001C_0004_002A_0016_0035_000D;
            @(posedge clkD) In_data = 256'h0036_0023_0035_002A_002D_000E_000B_0026_0041_0032_0030_002A_0015_001B_0007_0014;
            @(posedge clkD) In_data = 256'h0021_0020_0007_003B_003D_0022_0010_0023_002B_0023_0011_002B_0025_0023_0026_0018;
            @(posedge clkD) In_data = 256'h0022_003F_0017_002E_0011_0011_002B_002E_0031_002F_0030_0026_000A_0025_002B_0030;
            @(posedge clkD) In_data = 256'h0032_0021_0031_003F_001A_000C_000A_0001_0022_000E_001F_002B_0010_0040_002F_0000;
            @(posedge clkD) In_data = 256'h0036_0021_0030_0001_0015_0002_0032_0000_0026_0008_0038_003D_002D_0012_0019_000A;
            @(posedge clkD) In_data = 256'h0012_000B_0026_0024_0009_0002_001A_002E_000E_003A_0024_0013_0033_0029_0025_0007;
            @(posedge clkD) In_data = 256'h0023_000E_001B_001C_0035_0022_001A_0025_0001_003D_001F_0005_0015_0000_0024_0038;
            @(posedge clkD) In_data = 256'h0019_0021_0008_003E_0040_0022_0030_0025_0025_0005_003B_0018_0009_0007_002D_0006;
            @(posedge clkD) In_data = 256'h0032_003D_0036_0002_001B_0003_001E_002E_000C_0018_000F_0033_001B_0012_002F_0009;
            @(posedge clkD) In_data = 256'h003C_001D_0008_001B_0007_003D_0018_0025_0026_002F_003C_0018_0039_0016_0010_0004;
            @(posedge clkD) In_data = 256'h003F_0016_0014_0030_000E_000F_0003_002D_0000_0014_003A_002C_0028_0036_0011_0009;
            @(posedge clkD) In_data = 256'h0019_000B_002F_0011_0001_0014_0001_0019_0038_002E_0016_000F_002C_0021_0012_0009;
            @(posedge clkD) In_data = 256'h001E_0031_0022_0005_003A_0041_0005_0032_002B_0001_0029_000C_002E_0010_0001_002E;
            @(posedge clkD) In_data = 256'h002B_001A_0007_001D_0005_0041_0037_0000_000A_0041_003F_003E_0014_0027_0024_0000;
            @(posedge clkD) In_data = 256'h0001_0041_0034_002F_0020_002B_003C_0017_0003_0030_000A_003D_0010_0025_002C_003C;
            @(posedge clkD) In_data = 256'h0040_0006_002F_0040_0011_0000_0024_0024_001F_003E_0010_002B_001B_0000_0011_0025;
            @(posedge clkD) In_data = 256'h0013_000C_0009_0003_003E_0036_001B_0012_0039_0009_0002_0022_0002_0006_002D_0027;
            @(posedge clkD) In_data = 256'h0007_0018_0012_0030_0017_0008_0037_000C_0007_002D_001C_0002_0028_0039_0016_003F;
            @(posedge clkD) In_data = 256'h0034_0011_0035_002B_0003_0024_0003_0031_0028_0025_0005_0002_0013_002A_0037_003A;
            @(posedge clkD) In_data = 256'h0011_0001_002E_0029_001A_001D_0015_003F_002C_0040_0002_002F_0015_0036_000F_0007;
            @(posedge clkD) In_data = 256'h0015_000B_001A_003D_0040_001E_0034_003E_0006_0038_002F_0014_000B_001E_0007_0011;
            @(posedge clkD) In_data = 256'h0029_0034_0016_0022_0016_0006_002A_000B_0029_001A_0016_0005_002D_0028_002A_001A;
            @(posedge clkD) In_data = 256'h0003_001E_0003_0018_0004_0013_0014_003D_0038_0004_0004_000E_0041_0020_000C_0036;
            @(posedge clkD) In_data = 256'h0010_000E_0019_001B_000F_0003_003C_003B_0007_0002_000A_003A_003E_0008_0022_0025;
            @(posedge clkD) In_data = 256'h001B_002B_0010_0002_0010_0000_001D_000B_0029_0004_0027_0011_0022_003E_0004_0014;
            @(posedge clkD) In_data = 256'h003E_0030_003C_0017_0003_0007_002B_002B_0032_0022_0035_0010_0024_0019_0007_000B;
            @(posedge clkD) In_data = 256'h000E_0036_000D_0003_0036_0025_0003_002E_003D_001A_002B_0017_0023_002A_003A_002D;
            @(posedge clkD) In_data = 256'h0023_002E_003E_001A_001C_0040_0009_000A_001E_002B_001B_0005_0021_0029_001F_001E;
            @(posedge clkD) In_data = 256'h0041_0002_0020_000D_0014_002E_000D_0036_003C_0030_000E_002F_0022_0024_0009_002F;
            @(posedge clkD) In_data = 256'h001F_000A_0003_0032_0022_0004_0040_000A_0012_0036_0026_0009_0016_001C_0029_0010;
            @(posedge clkD) In_data = 256'h003D_0034_0009_0026_002B_0030_003D_0007_0011_0019_0037_0040_0037_0038_0026_002C;
            @(posedge clkD) In_data = 256'h0024_0040_002C_003D_003E_003E_0020_0023_0011_002A_0017_003C_002C_001D_0034_000D;
            @(posedge clkD) In_data = 256'h0033_0038_003A_0019_0012_0038_0008_0010_003A_0009_0022_001C_003F_002F_000A_0014;
            @(posedge clkD) In_data = 256'h0035_001E_0025_0022_002C_0037_0021_0008_001C_0005_0030_0010_002B_0023_002F_0016;
            @(posedge clkD) In_data = 256'h001E_002D_0027_0023_0034_0006_001E_0025_002F_0022_0028_0026_0018_002B_0034_003C;
            @(posedge clkD) In_data = 256'h0014_002A_0014_0006_0013_0030_002B_0025_0028_0010_002E_003B_0010_000A_0019_000A;
            @(posedge clkD) In_data = 256'h0037_002F_0006_0013_0021_0036_0003_0019_001A_0011_0005_003B_0036_0002_0037_0002;
            @(posedge clkD) In_data = 256'h0002_0000_001D_0007_000D_0002_0015_0008_0030_003B_001B_0028_0022_003D_0031_0030;
            @(posedge clkD) In_data = 256'h0006_0032_0026_003D_0034_0001_0008_001D_0034_000E_0029_0034_0041_0014_0017_0037;
            @(posedge clkD) In_data = 256'h0038_0027_0035_0019_0032_0011_0034_0024_003C_0016_000A_0015_0003_0038_0015_0017;
            @(posedge clkD) In_data = 256'h0005_0041_0004_003F_0005_003F_0026_0013_002D_001E_0038_0010_0015_0037_0027_0031;
            @(posedge clkD) In_data = 256'h0005_003C_003C_0027_0027_0016_0005_0032_002A_0009_0003_001A_0015_001F_0005_0009;
            @(posedge clkD) In_data = 256'h0005_0040_0013_0032_002B_000D_0034_000F_0000_000E_0007_0013_0037_002F_002C_0027;
            @(posedge clkD) In_data = 256'h003C_0025_002C_000F_0028_003D_0010_003E_0021_002E_001F_0006_0039_002D_0011_0020;
            @(posedge clkD) In_data = 256'h0039_0030_000E_0020_0004_0033_003B_0002_0000_0000_0000_0000_0000_0000_0000_0000;
        end   
        // end of packet
        // @(posedge clkD)
        //output is ready
        

        // @(posedge clkD) Out_ready   =   1'b1 ;
         
        // while (!In_ready)  


            // 9th

        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;

                            In_data = 256'h0006_0035_0017_0015_0003_001B_002E_0020_0004_003C_0017_0010_0014_0023_0026_000C ;
            @(posedge clkD) In_data = 256'h0036_0010_0007_0015_003F_0002_000C_0016_0002_000C_0000_003B_0037_003E_0021_0040 ;
            @(posedge clkD) In_data = 256'h0000_0041_0003_0002_0034_0037_003E_000D_0030_000B_0004_0016_0020_001C_0034_0007 ;
            @(posedge clkD) In_data = 256'h000E_002F_0014_0032_001E_0041_000E_000A_000F_0019_0002_000E_0024_0037_0040_0035 ;
            @(posedge clkD) In_data = 256'h0002_003B_0041_002F_0029_0038_0015_0036_0020_000F_0011_001D_000E_0007_0030_003B ;
            @(posedge clkD) In_data = 256'h0040_0025_0030_0005_0041_0011_0005_002D_0020_0031_0023_003A_0023_0007_0005_003C ;
            @(posedge clkD) In_data = 256'h0031_0036_001C_0001_0015_0010_0007_0034_002A_000E_0030_0025_000F_0039_000C_0039 ;
            @(posedge clkD) In_data = 256'h0008_0007_002C_0005_0001_0006_0035_0028_000F_000A_003E_0001_001E_0017_0019_0014 ;
            @(posedge clkD) In_data = 256'h000C_0036_000C_0038_0017_002A_003B_0019_003E_002B_001F_003B_0004_0020_003D_002B ;
            @(posedge clkD) In_data = 256'h0021_002B_003E_0011_0006_0037_0022_0026_001C_0006_0034_0028_003A_0035_0041_0014 ;
            @(posedge clkD) In_data = 256'h003E_0029_0035_0013_003C_003E_0011_003D_003A_0035_0033_0008_0010_002F_0013_0009 ;
            @(posedge clkD) In_data = 256'h0022_002B_0011_0026_0002_003C_0032_001D_0015_002C_0036_0017_0012_0028_0034_0016 ;
            @(posedge clkD) In_data = 256'h001A_0034_003F_0022_0032_0038_000B_000D_0001_002E_000D_0036_0018_0002_0025_0013 ;
            @(posedge clkD) In_data = 256'h0033_000C_003F_003A_000F_0023_0008_0002_0009_0018_0011_0006_0018_0012_0000_0011 ;
            @(posedge clkD) In_data = 256'h0035_0014_000F_001E_000F_0007_0012_0023_0008_0031_001A_0004_0041_0013_0016_001C ;
            @(posedge clkD) In_data = 256'h0006_000E_0022_0006_0016_0010_0018_000F_0024_0007_0003_001B_003F_003A_001C_0002 ;
            @(posedge clkD) In_data = 256'h001C_0013_0030_0004_0040_002C_0009_0028_000B_0037_0031_003C_003E_0023_0029_0006 ;
            @(posedge clkD) In_data = 256'h0008_0026_001A_0014_002F_002C_0006_0041_001B_0013_0020_0019_0031_001F_0038_000E ;
            @(posedge clkD) In_data = 256'h0025_003C_0039_0011_0032_003B_0039_001D_0021_001F_0017_000A_000D_001F_002A_0034 ;
            @(posedge clkD) In_data = 256'h0009_0009_0041_003F_000D_003E_0032_002C_001F_001C_0011_0006_0022_001C_0006_000D ;
            @(posedge clkD) In_data = 256'h0031_0023_001F_000C_0029_002C_000B_0037_003C_002B_0030_0016_003A_000F_000E_0005 ;
            @(posedge clkD) In_data = 256'h0019_0037_003C_001E_0039_0026_0016_003E_0035_001C_002A_0000_0017_000E_002B_0006 ;
            @(posedge clkD) In_data = 256'h001D_0033_0020_000C_0015_001A_0037_003A_0028_001F_002E_001D_0001_0005_0022_003E ;
            @(posedge clkD) In_data = 256'h0022_000D_0022_003D_0005_0001_0023_0038_001E_0040_0034_003C_001C_0026_002D_0010 ;
            @(posedge clkD) In_data = 256'h0036_002A_003B_000D_000A_001D_000F_003C_0038_003E_0010_0011_0023_0002_003A_003D ;
            @(posedge clkD) In_data = 256'h0034_0034_0036_0020_0030_0014_0011_0031_0035_0017_0019_0038_003D_003C_0036_000F ;
            @(posedge clkD) In_data = 256'h002A_0008_002B_0040_0026_0017_0034_0004_0009_0021_001E_0002_002C_003F_003A_000E ;
            @(posedge clkD) In_data = 256'h0027_0040_001F_0002_0019_0027_000D_0024_002C_000B_003F_002E_0022_0000_0030_000D ;
            @(posedge clkD) In_data = 256'h001D_0021_0008_0011_000C_002C_0037_0032_0010_002D_0007_000A_0004_0003_001F_0033 ;
            @(posedge clkD) In_data = 256'h002D_0028_0023_000B_0001_0011_0006_003E_0039_0026_0012_0018_0028_000A_0002_0029 ;
            @(posedge clkD) In_data = 256'h0015_0021_0011_000B_003B_0039_0021_001C_001C_000A_0024_003D_0021_000B_003D_001B ;
            @(posedge clkD) In_data = 256'h003B_000D_001A_0026_003E_000D_002C_0007_000C_0039_0019_0008_0039_0006_0033_002D ;
            @(posedge clkD) In_data = 256'h0040_0026_0020_0035_000F_002B_0018_0040_0033_000F_0021_002E_0029_0013_0041_0021 ;
            @(posedge clkD) In_data = 256'h0020_0020_0000_0035_0014_003C_0008_0029_0023_0007_0028_0003_001B_0041_003B_0017 ;
            @(posedge clkD) In_data = 256'h0030_0037_0002_001D_0012_0015_003F_001D_0011_0015_0033_0012_0012_0002_0012_000A ;
            @(posedge clkD) In_data = 256'h002C_002A_0015_0031_0016_000D_0025_0022_0037_0008_0023_000C_0034_0032_0040_0003 ;
            @(posedge clkD) In_data = 256'h000C_001B_0041_0025_002F_0032_003D_0004_0022_0010_003B_0035_0002_0031_0021_0032 ;
            @(posedge clkD) In_data = 256'h003A_0007_0023_0014_003A_0002_001F_003D_001A_000B_000C_0025_0011_0024_0041_002F ;
            @(posedge clkD) In_data = 256'h0026_002D_001D_0028_0001_001F_0037_003E_002E_0022_0033_0021_0039_0040_0007_0033 ;
            @(posedge clkD) In_data = 256'h001B_0017_0031_0008_0029_0015_0008_0003_0024_0034_002F_000F_003F_001F_002C_0004 ;
            @(posedge clkD) In_data = 256'h0040_0014_000B_0014_000C_003B_0007_0010_0031_0012_0004_002B_0032_001A_001C_003E ;
            @(posedge clkD) In_data = 256'h0000_0012_002B_0006_0003_0014_0014_003E_0025_000E_0012_001B_000B_003B_0031_0000 ;
            @(posedge clkD) In_data = 256'h0027_003B_001F_000A_0001_0024_002B_0013_0027_000F_0037_003D_003D_0028_000A_001F ;
            @(posedge clkD) In_data = 256'h001C_0033_0037_0023_001F_0022_0032_001B_0018_0030_0022_0003_0022_0015_000E_0040 ;
            @(posedge clkD) In_data = 256'h0022_0028_0026_0022_0006_0006_000F_000D_0028_0022_0013_0031_0025_0036_001C_001A ;
            @(posedge clkD) In_data = 256'h001A_000F_0021_000A_0018_001D_0036_001B_0039_0035_0026_000C_0006_0029_000D_0011 ;
            @(posedge clkD) In_data = 256'h0022_001E_001F_000C_0025_0020_0031_0029_003E_001A_002B_0010_003B_0017_0025_001C ;
            @(posedge clkD) In_data = 256'h000E_0023_0014_0033_0017_0000_0002_003C_003C_001E_0014_0015_0010_0012_001D_0039 ;
            @(posedge clkD) In_data = 256'h0001_003E_003B_0037_0003_003C_0021_003E_0037_0037_0031_0040_001A_0035_000B_0032 ;
            @(posedge clkD) In_data = 256'h002F_0032_0017_001E_0005_003E_0011_0012_0030_000C_003B_003B_0003_0019_003E_0031 ;
            @(posedge clkD) In_data = 256'h0022_0006_0017_0036_003C_0014_0041_0030_0025_001D_0037_0036_003A_001D_000D_0035 ;
            @(posedge clkD) In_data = 256'h002B_000C_001E_0007_001D_0017_0032_003D_0002_0018_003F_0016_000E_0009_002D_000B ;
            @(posedge clkD) In_data = 256'h0028_001D_0023_0004_0025_001C_000C_0016_000D_0039_003F_0028_0017_001B_0007_0018 ;
            @(posedge clkD) In_data = 256'h0033_001E_0011_002F_0032_0021_000A_0038_000A_001E_0006_0039_0002_0023_0000_0041 ;
            @(posedge clkD) In_data = 256'h0003_001A_0029_0029_0005_0007_000A_001B_002E_0029_0026_0030_0029_003D_002E_000D ;
            @(posedge clkD) In_data = 256'h000B_0037_0000_0021_001B_0010_003B_0020_001E_001A_0024_0037_000D_0024_0027_0037 ;
            @(posedge clkD) In_data = 256'h0002_0002_0016_0002_0009_0018_000D_0010_0027_001C_0031_0021_0006_003B_000B_0036 ;
            @(posedge clkD) In_data = 256'h002B_001C_0005_0040_002B_0023_0009_0035_003C_003E_002F_0013_003B_002A_0014_0040 ;
            @(posedge clkD) In_data = 256'h0018_0035_003A_000E_0040_0024_0010_0028_0035_0000_0021_0025_0030_0028_000F_0002 ;
            @(posedge clkD) In_data = 256'h0012_001F_0033_003D_002F_003D_0014_003D_0016_000B_0036_002A_0012_001A_000D_002A ;
            @(posedge clkD) In_data = 256'h0028_0014_000D_0020_0033_002D_0005_0024_0040_001F_0029_0001_0020_001A_0028_0016 ;
            @(posedge clkD) In_data = 256'h0027_002F_0014_002C_002B_0005_0003_0039_003F_0007_002C_002C_0002_003A_0033_0037 ;
            @(posedge clkD) In_data = 256'h0041_0014_0012_0040_0021_001D_0037_0023_0000_0000_0000_0000_0000_0000_0000_0000 ;
            
       
       
       
       
       



       


        end

        if (In_ready) begin
            @(posedge clkD) In_valid    <=      1'b1;
                            In_data = 256'h0010_003C_000F_002B_0010_000D_0016_000A_000E_0028_002D_0013_002B_0028_001E_0025;
            @(posedge clkD) In_data = 256'h001B_001F_0032_0008_003A_0002_000C_0035_0027_0011_0033_0021_0033_003D_002B_0025;
            @(posedge clkD) In_data = 256'h0002_0004_0006_0007_0041_0006_0014_0009_000C_0004_0015_0013_0037_0020_000B_0032;
            @(posedge clkD) In_data = 256'h001A_0015_0039_0023_0012_0032_0013_0037_000F_0011_0003_003C_0041_0032_002D_0016;
            @(posedge clkD) In_data = 256'h0041_003D_0025_0039_002A_001B_002C_0011_0020_0005_0013_0005_002D_0019_0038_0001;
            @(posedge clkD) In_data = 256'h000A_0024_000B_002E_002A_003B_002B_000A_0000_000D_0004_003A_0012_0019_0020_001F;
            @(posedge clkD) In_data = 256'h0022_003F_003F_0018_003F_002D_003F_0024_0024_0004_0026_003B_0024_0037_001A_000F;
            @(posedge clkD) In_data = 256'h0015_0027_0000_0029_003F_003F_000A_002E_003D_0033_0003_0027_0009_0006_0017_0013;
            @(posedge clkD) In_data = 256'h000D_002D_000F_0024_0039_0039_003E_0025_002C_0000_000F_001B_000A_0036_002E_0032;
            @(posedge clkD) In_data = 256'h0027_0034_0007_0017_0018_003E_000A_0039_0024_003A_0005_0016_003F_0034_0028_0031;
            @(posedge clkD) In_data = 256'h001F_0001_0017_002F_0025_003D_0016_0027_0017_001B_000E_0011_002D_0034_0013_003A;
            @(posedge clkD) In_data = 256'h0009_0013_003B_0017_0035_0001_0030_0007_0040_0017_002D_0011_003D_0001_0007_003B;
            @(posedge clkD) In_data = 256'h0015_0033_000B_000E_0024_0032_003F_0041_003F_000E_0003_0033_0013_0001_0025_0006;
            @(posedge clkD) In_data = 256'h0016_0034_0000_003C_002C_0000_0035_002F_002C_003F_0027_0017_0029_0031_003F_0028;
            @(posedge clkD) In_data = 256'h0025_000E_002D_001F_000D_001F_000B_001C_0019_0009_0018_0032_0019_0009_000D_0033;
            @(posedge clkD) In_data = 256'h0007_0039_003F_0002_0019_0031_002B_0028_0010_0023_0002_0008_002F_003D_0030_0009;
            @(posedge clkD) In_data = 256'h0035_001F_002D_0036_0037_001D_0033_0022_0038_0041_002D_000F_0037_0032_0017_0041;
            @(posedge clkD) In_data = 256'h0038_0009_002E_0001_0012_0015_0014_0029_001F_001D_0013_0027_000F_0032_0033_0008;
            @(posedge clkD) In_data = 256'h001D_0023_0041_001F_0021_0020_0031_002F_0027_0033_002C_0035_000C_0001_0034_0012;
            @(posedge clkD) In_data = 256'h002C_0024_000A_0007_0016_000D_0039_001B_0032_001A_003E_000C_0013_0037_002F_0028;
            @(posedge clkD) In_data = 256'h000C_001A_002B_0034_0019_0027_0007_000E_0031_001F_003C_0017_000B_000F_0000_0036;
            @(posedge clkD) In_data = 256'h0038_0006_000A_0007_0017_002C_002A_0004_0026_0033_0030_0021_0003_0036_003A_001B;
            @(posedge clkD) In_data = 256'h001F_0024_0038_0020_001C_0034_003C_0028_0033_0035_001B_0011_0019_0026_0024_001F;
            @(posedge clkD) In_data = 256'h0011_003B_0028_001C_003B_0035_0011_0016_0022_0009_0008_0027_0021_0018_001A_0038;
            @(posedge clkD) In_data = 256'h003F_001B_0015_0041_002B_000C_0017_001C_0018_0040_0001_000C_0005_0030_0022_002E;
            @(posedge clkD) In_data = 256'h001D_003B_002B_0040_0024_001B_002B_0035_0026_000F_000D_000C_0035_0022_0041_0008;
            @(posedge clkD) In_data = 256'h0021_0038_0020_0034_0014_000D_002C_0011_000E_003E_003C_0014_0013_001C_000B_000A;
            @(posedge clkD) In_data = 256'h001E_003E_0006_0033_003C_0007_0008_0017_003D_000B_0020_0005_0000_0028_0012_000A;
            @(posedge clkD) In_data = 256'h0002_000E_000E_0027_003A_0012_002F_003E_0038_0026_000E_003E_0009_0003_003A_002E;
            @(posedge clkD) In_data = 256'h0039_0007_002A_0029_003F_0012_002C_0014_002E_0023_002F_0013_0030_001E_0014_001F;
            @(posedge clkD) In_data = 256'h0029_0009_0011_0020_002F_0040_0034_0038_002D_0013_0007_0016_0010_0013_003C_0005;
            @(posedge clkD) In_data = 256'h0027_0006_0001_000F_0034_0009_001A_002E_0019_0001_0006_0029_0001_0005_0004_0012;
            @(posedge clkD) In_data = 256'h001D_002D_003F_0015_000F_000C_001F_0026_0016_0015_0020_0027_0030_0035_001A_0016;
            @(posedge clkD) In_data = 256'h0027_002F_0036_0023_0029_0034_0031_0033_0005_0022_0026_0020_0011_0032_0005_0020;
            @(posedge clkD) In_data = 256'h0029_0033_002C_0016_0032_0030_0018_002A_0036_0000_000B_0020_0039_0011_0003_0012;
            @(posedge clkD) In_data = 256'h003D_0013_002B_0035_0019_000E_0028_0014_000D_001E_0014_0024_0007_0004_000B_0028;
            @(posedge clkD) In_data = 256'h001B_0000_0022_0023_0013_0008_0003_0005_0036_0027_003D_000E_0031_0022_0039_0024;
            @(posedge clkD) In_data = 256'h0004_000A_0032_0017_003B_0039_001A_0015_0025_000C_0005_000C_0016_0030_0024_001A;
            @(posedge clkD) In_data = 256'h0037_000D_001B_0009_0006_0008_0032_0015_0015_0016_0031_0008_0036_0019_0031_0029;
            @(posedge clkD) In_data = 256'h0002_0011_0005_003A_0016_0025_003F_0041_0038_003F_000A_001A_0034_003E_003E_0020;
            @(posedge clkD) In_data = 256'h0010_0000_002D_0028_0023_003A_0016_0006_000C_0009_0004_0035_0002_0032_0000_0041;
            @(posedge clkD) In_data = 256'h003B_0019_002F_000D_0006_0041_0011_002D_0000_0001_000E_0018_003F_0024_000D_002C;
            @(posedge clkD) In_data = 256'h0040_0026_0006_0031_003D_001E_0007_0018_0038_003E_002B_0040_0016_001C_001B_001D;
            @(posedge clkD) In_data = 256'h003D_0033_0031_0029_0038_0028_0033_0014_0021_002B_0006_0023_0036_0033_0028_001D;
            @(posedge clkD) In_data = 256'h0041_001D_0038_0003_003E_0019_000D_001F_0033_0003_000D_0032_0028_003D_0007_0010;
            @(posedge clkD) In_data = 256'h003B_001D_003B_0039_0015_0023_001B_003B_0033_0018_003A_001A_001D_0010_0011_0036;
            @(posedge clkD) In_data = 256'h0021_003C_0012_0012_0026_0020_002D_0024_0020_0004_001B_0019_002C_003F_0007_001F;
            @(posedge clkD) In_data = 256'h0017_0040_0017_0034_003A_000A_0024_0033_0036_002B_0022_0031_002A_0001_002B_0007;
            @(posedge clkD) In_data = 256'h0021_0011_0005_0032_0029_0032_000D_0005_0001_0011_0002_0020_003D_0025_001F_001E;
            @(posedge clkD) In_data = 256'h002F_000D_002A_002F_0036_0013_002D_0020_0041_003C_000F_0003_001D_0012_0034_0011;
            @(posedge clkD) In_data = 256'h0038_0020_0017_001D_003A_0033_0039_0015_001B_0015_0031_0026_002B_001C_0020_0025;
            @(posedge clkD) In_data = 256'h000C_001F_0030_0022_0025_0022_0020_003F_0021_0005_0038_003D_0021_0001_0023_0013;
            @(posedge clkD) In_data = 256'h0016_0010_003B_003E_0016_0033_0018_003E_001C_000E_002B_002B_002B_002A_0009_000C;
            @(posedge clkD) In_data = 256'h0034_002C_0001_003D_0002_0006_0030_000B_0006_0004_000A_0036_003F_0030_002C_0030;
            @(posedge clkD) In_data = 256'h0037_001A_001A_002B_0033_002C_0004_0040_0008_0006_003E_002F_003C_0035_002E_000D;
            @(posedge clkD) In_data = 256'h0009_0003_0003_0022_0024_0021_0004_0020_0026_001F_0019_0007_003C_0033_0017_0027;
            @(posedge clkD) In_data = 256'h0024_0035_0032_0033_0026_000E_0015_000E_0029_0004_0022_001E_0020_0029_0027_0021;
            @(posedge clkD) In_data = 256'h0024_002B_0010_0008_0026_0008_003F_0026_001D_0012_0012_0032_003F_002E_000A_0029;
            @(posedge clkD) In_data = 256'h0029_0019_0037_0030_0031_000F_001C_0009_001C_003D_0008_0009_0002_0004_0033_0040;
            @(posedge clkD) In_data = 256'h0015_001B_0022_002D_0019_000F_002D_0032_001A_0033_0026_0037_0039_000E_0024_000E;
            @(posedge clkD) In_data = 256'h002F_000E_0024_0019_0027_0041_0026_003A_0040_000A_001E_003F_001C_001E_002A_003F;
            @(posedge clkD) In_data = 256'h0011_000B_002A_0034_0011_002C_0021_0018_0016_002D_0015_0017_003D_0036_000D_002C;
            @(posedge clkD) In_data = 256'h0037_0040_0007_0018_0032_001E_003A_0020_0000_0000_0000_0000_0000_0000_0000_0000;
        end   


        @(posedge clkD) In_valid    <=      1'b1;
        
        @(posedge clkD) In_valid    <=      1'b1;
        Out_ready   =   1'b1 ; 
        while (!In_ready)    ;
        #3000 $finish();   
     
     end 
    
endmodule